<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-29.6556,3.8211,53.5444,-88.5789</PageViewport>
<gate>
<ID>2</ID>
<type>AA_INVERTER</type>
<position>15,-9</position>
<input>
<ID>IN_0</ID>1 </input>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>4,-9</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>-2,-17</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>7</ID>
<type>AA_INVERTER</type>
<position>15,-17</position>
<input>
<ID>IN_0</ID>2 </input>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>9</ID>
<type>AA_AND2</type>
<position>28.5,-10</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>17 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>11</ID>
<type>AA_AND2</type>
<position>28.5,-16</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>18 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>31</ID>
<type>BE_NOR2</type>
<position>42.5,-12.5</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>18 </input>
<output>
<ID>OUT</ID>37 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>32</ID>
<type>AA_INVERTER</type>
<position>15,-25.5</position>
<input>
<ID>IN_0</ID>19 </input>
<output>
<ID>OUT_0</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>33</ID>
<type>AA_TOGGLE</type>
<position>4,-25.5</position>
<output>
<ID>OUT_0</ID>19 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>34</ID>
<type>AA_TOGGLE</type>
<position>-2,-33.5</position>
<output>
<ID>OUT_0</ID>20 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>35</ID>
<type>AA_INVERTER</type>
<position>15,-33.5</position>
<input>
<ID>IN_0</ID>20 </input>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>36</ID>
<type>AA_AND2</type>
<position>28.5,-26.5</position>
<input>
<ID>IN_0</ID>22 </input>
<input>
<ID>IN_1</ID>20 </input>
<output>
<ID>OUT</ID>23 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>37</ID>
<type>AA_AND2</type>
<position>28.5,-32.5</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>24 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>38</ID>
<type>BE_NOR2</type>
<position>42.5,-29</position>
<input>
<ID>IN_0</ID>23 </input>
<input>
<ID>IN_1</ID>24 </input>
<output>
<ID>OUT</ID>38 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>39</ID>
<type>AA_INVERTER</type>
<position>15,-43</position>
<input>
<ID>IN_0</ID>25 </input>
<output>
<ID>OUT_0</ID>28 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>40</ID>
<type>AA_TOGGLE</type>
<position>4,-43</position>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>41</ID>
<type>AA_TOGGLE</type>
<position>-2,-50.5</position>
<output>
<ID>OUT_0</ID>26 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>42</ID>
<type>AA_INVERTER</type>
<position>15,-51</position>
<input>
<ID>IN_0</ID>26 </input>
<output>
<ID>OUT_0</ID>27 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>43</ID>
<type>AA_AND2</type>
<position>28.5,-44</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>29 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_AND2</type>
<position>28.5,-50</position>
<input>
<ID>IN_0</ID>25 </input>
<input>
<ID>IN_1</ID>27 </input>
<output>
<ID>OUT</ID>30 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>45</ID>
<type>BE_NOR2</type>
<position>42.5,-46.5</position>
<input>
<ID>IN_0</ID>29 </input>
<input>
<ID>IN_1</ID>30 </input>
<output>
<ID>OUT</ID>40 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>46</ID>
<type>AA_INVERTER</type>
<position>15.5,-60.5</position>
<input>
<ID>IN_0</ID>31 </input>
<output>
<ID>OUT_0</ID>34 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>47</ID>
<type>AA_TOGGLE</type>
<position>4.5,-60.5</position>
<output>
<ID>OUT_0</ID>31 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>48</ID>
<type>AA_TOGGLE</type>
<position>-1.5,-69</position>
<output>
<ID>OUT_0</ID>32 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>49</ID>
<type>AA_INVERTER</type>
<position>15.5,-68.5</position>
<input>
<ID>IN_0</ID>32 </input>
<output>
<ID>OUT_0</ID>33 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>50</ID>
<type>AA_AND2</type>
<position>29,-61.5</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_1</ID>32 </input>
<output>
<ID>OUT</ID>35 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>51</ID>
<type>AA_AND2</type>
<position>29,-67.5</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>33 </input>
<output>
<ID>OUT</ID>36 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>52</ID>
<type>BE_NOR2</type>
<position>43,-64.5</position>
<input>
<ID>IN_0</ID>35 </input>
<input>
<ID>IN_1</ID>36 </input>
<output>
<ID>OUT</ID>42 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>54</ID>
<type>AA_AND2</type>
<position>59.5,-24.5</position>
<input>
<ID>IN_0</ID>37 </input>
<input>
<ID>IN_1</ID>23 </input>
<output>
<ID>OUT</ID>50 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>56</ID>
<type>AA_AND2</type>
<position>59.5,-36</position>
<input>
<ID>IN_0</ID>37 </input>
<input>
<ID>IN_1</ID>24 </input>
<output>
<ID>OUT</ID>46 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>64</ID>
<type>AA_AND3</type>
<position>59.5,-42.5</position>
<input>
<ID>IN_0</ID>37 </input>
<input>
<ID>IN_1</ID>38 </input>
<input>
<ID>IN_2</ID>29 </input>
<output>
<ID>OUT</ID>49 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>66</ID>
<type>AA_AND3</type>
<position>59.5,-52</position>
<input>
<ID>IN_0</ID>37 </input>
<input>
<ID>IN_1</ID>38 </input>
<input>
<ID>IN_2</ID>30 </input>
<output>
<ID>OUT</ID>45 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>68</ID>
<type>AA_AND4</type>
<position>59.5,-59.5</position>
<input>
<ID>IN_0</ID>37 </input>
<input>
<ID>IN_1</ID>38 </input>
<input>
<ID>IN_2</ID>40 </input>
<input>
<ID>IN_3</ID>35 </input>
<output>
<ID>OUT</ID>48 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>70</ID>
<type>AA_AND4</type>
<position>59.5,-70</position>
<input>
<ID>IN_0</ID>37 </input>
<input>
<ID>IN_1</ID>38 </input>
<input>
<ID>IN_2</ID>40 </input>
<input>
<ID>IN_3</ID>36 </input>
<output>
<ID>OUT</ID>44 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>72</ID>
<type>AA_AND4</type>
<position>59.5,-79</position>
<input>
<ID>IN_0</ID>37 </input>
<input>
<ID>IN_1</ID>38 </input>
<input>
<ID>IN_2</ID>40 </input>
<input>
<ID>IN_3</ID>42 </input>
<output>
<ID>OUT</ID>43 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>74</ID>
<type>AE_OR4</type>
<position>80,-34.5</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>50 </input>
<input>
<ID>IN_2</ID>49 </input>
<input>
<ID>IN_3</ID>48 </input>
<output>
<ID>OUT</ID>51 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>76</ID>
<type>AE_OR4</type>
<position>80,-51</position>
<input>
<ID>IN_0</ID>18 </input>
<input>
<ID>IN_1</ID>46 </input>
<input>
<ID>IN_2</ID>45 </input>
<input>
<ID>IN_3</ID>44 </input>
<output>
<ID>OUT</ID>47 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>78</ID>
<type>GA_LED</type>
<position>89,-36</position>
<input>
<ID>N_in0</ID>51 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>82</ID>
<type>GA_LED</type>
<position>89,-51.5</position>
<input>
<ID>N_in0</ID>47 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>84</ID>
<type>GA_LED</type>
<position>89,-78.5</position>
<input>
<ID>N_in0</ID>43 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>86</ID>
<type>AA_LABEL</type>
<position>-1,-8.5</position>
<gparam>LABEL_TEXT A3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>87</ID>
<type>AA_LABEL</type>
<position>-7,-16.5</position>
<gparam>LABEL_TEXT B3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>88</ID>
<type>AA_LABEL</type>
<position>0,-25.5</position>
<gparam>LABEL_TEXT A2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>89</ID>
<type>AA_LABEL</type>
<position>-7.5,-33</position>
<gparam>LABEL_TEXT B2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>90</ID>
<type>AA_LABEL</type>
<position>0,-42.5</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>91</ID>
<type>AA_LABEL</type>
<position>-7,-50</position>
<gparam>LABEL_TEXT B1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>92</ID>
<type>AA_LABEL</type>
<position>0.5,-60</position>
<gparam>LABEL_TEXT A0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>93</ID>
<type>AA_LABEL</type>
<position>-6.5,-68.5</position>
<gparam>LABEL_TEXT B0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>95</ID>
<type>AA_LABEL</type>
<position>99.5,-35.5</position>
<gparam>LABEL_TEXT AB</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>97</ID>
<type>AA_LABEL</type>
<position>100,-51</position>
<gparam>LABEL_TEXT A>B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>99</ID>
<type>AA_LABEL</type>
<position>99,-78</position>
<gparam>LABEL_TEXT A=B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>6,-9,12,-9</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>9 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>9,-12.5,9,-9</points>
<intersection>-12.5 7</intersection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>9,-12.5,25.5,-12.5</points>
<intersection>9 6</intersection>
<intersection>25.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>25.5,-15,25.5,-12.5</points>
<connection>
<GID>11</GID>
<name>IN_0</name></connection>
<intersection>-12.5 7</intersection></vsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>0,-17,12,-17</points>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>9 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>9,-17,9,-13.5</points>
<intersection>-17 1</intersection>
<intersection>-13.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>9,-13.5,24,-13.5</points>
<intersection>9 6</intersection>
<intersection>24 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>24,-13.5,24,-11</points>
<intersection>-13.5 7</intersection>
<intersection>-11 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>24,-11,25.5,-11</points>
<connection>
<GID>9</GID>
<name>IN_1</name></connection>
<intersection>24 8</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>18,-17,25.5,-17</points>
<connection>
<GID>11</GID>
<name>IN_1</name></connection>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>18,-9,25.5,-9</points>
<connection>
<GID>9</GID>
<name>IN_0</name></connection>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-10,35.5,-7</points>
<intersection>-10 2</intersection>
<intersection>-7 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35.5,-7,77,-7</points>
<intersection>35.5 0</intersection>
<intersection>39.5 4</intersection>
<intersection>77 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>31.5,-10,35.5,-10</points>
<connection>
<GID>9</GID>
<name>OUT</name></connection>
<intersection>35.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>77,-31.5,77,-7</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<intersection>-7 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>39.5,-11.5,39.5,-7</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>-7 1</intersection></vsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-19,35.5,-16</points>
<intersection>-19 1</intersection>
<intersection>-16 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35.5,-19,69,-19</points>
<intersection>35.5 0</intersection>
<intersection>39.5 5</intersection>
<intersection>69 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>31.5,-16,35.5,-16</points>
<connection>
<GID>11</GID>
<name>OUT</name></connection>
<intersection>35.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>69,-48,69,-19</points>
<intersection>-48 4</intersection>
<intersection>-19 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>69,-48,77,-48</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<intersection>69 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>39.5,-19,39.5,-13.5</points>
<connection>
<GID>31</GID>
<name>IN_1</name></connection>
<intersection>-19 1</intersection></vsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>6,-25.5,12,-25.5</points>
<connection>
<GID>33</GID>
<name>OUT_0</name></connection>
<connection>
<GID>32</GID>
<name>IN_0</name></connection>
<intersection>8.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>8.5,-29,8.5,-25.5</points>
<intersection>-29 7</intersection>
<intersection>-25.5 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>8.5,-29,25,-29</points>
<intersection>8.5 6</intersection>
<intersection>25 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>25,-31.5,25,-29</points>
<intersection>-31.5 11</intersection>
<intersection>-29 7</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>25,-31.5,25.5,-31.5</points>
<connection>
<GID>37</GID>
<name>IN_0</name></connection>
<intersection>25 8</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>0,-33.5,12,-33.5</points>
<connection>
<GID>35</GID>
<name>IN_0</name></connection>
<connection>
<GID>34</GID>
<name>OUT_0</name></connection>
<intersection>9 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>9,-33.5,9,-30</points>
<intersection>-33.5 1</intersection>
<intersection>-30 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>9,-30,24,-30</points>
<intersection>9 6</intersection>
<intersection>24 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>24,-30,24,-27.5</points>
<intersection>-30 7</intersection>
<intersection>-27.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>24,-27.5,25.5,-27.5</points>
<connection>
<GID>36</GID>
<name>IN_1</name></connection>
<intersection>24 8</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>18,-33.5,25.5,-33.5</points>
<connection>
<GID>35</GID>
<name>OUT_0</name></connection>
<connection>
<GID>37</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>18,-25.5,25.5,-25.5</points>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection>
<connection>
<GID>36</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-26.5,35.5,-25.5</points>
<intersection>-26.5 2</intersection>
<intersection>-25.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35.5,-25.5,56.5,-25.5</points>
<connection>
<GID>54</GID>
<name>IN_1</name></connection>
<intersection>35.5 0</intersection>
<intersection>38.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>31.5,-26.5,35.5,-26.5</points>
<connection>
<GID>36</GID>
<name>OUT</name></connection>
<intersection>35.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>38.5,-28,38.5,-25.5</points>
<intersection>-28 5</intersection>
<intersection>-25.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>38.5,-28,39.5,-28</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>38.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-37,35.5,-30</points>
<intersection>-37 1</intersection>
<intersection>-32.5 2</intersection>
<intersection>-30 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35.5,-37,56.5,-37</points>
<connection>
<GID>56</GID>
<name>IN_1</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>31.5,-32.5,35.5,-32.5</points>
<connection>
<GID>37</GID>
<name>OUT</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>35.5,-30,39.5,-30</points>
<connection>
<GID>38</GID>
<name>IN_1</name></connection>
<intersection>35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>6,-43,12,-43</points>
<connection>
<GID>40</GID>
<name>OUT_0</name></connection>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>9 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>9,-46.5,9,-43</points>
<intersection>-46.5 7</intersection>
<intersection>-43 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>9,-46.5,25.5,-46.5</points>
<intersection>9 6</intersection>
<intersection>25.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>25.5,-49,25.5,-46.5</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>-46.5 7</intersection></vsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>0,-50.5,12,-50.5</points>
<connection>
<GID>41</GID>
<name>OUT_0</name></connection>
<intersection>9 6</intersection>
<intersection>12 12</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>9,-50.5,9,-47.5</points>
<intersection>-50.5 1</intersection>
<intersection>-47.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>9,-47.5,24,-47.5</points>
<intersection>9 6</intersection>
<intersection>24 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>24,-47.5,24,-45</points>
<intersection>-47.5 7</intersection>
<intersection>-45 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>24,-45,25.5,-45</points>
<connection>
<GID>43</GID>
<name>IN_1</name></connection>
<intersection>24 8</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>12,-51,12,-50.5</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>-50.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>18,-51,25.5,-51</points>
<connection>
<GID>44</GID>
<name>IN_1</name></connection>
<connection>
<GID>42</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>18,-43,25.5,-43</points>
<connection>
<GID>43</GID>
<name>IN_0</name></connection>
<connection>
<GID>39</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-45.5,35.5,-43.5</points>
<intersection>-45.5 5</intersection>
<intersection>-44 2</intersection>
<intersection>-43.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35.5,-43.5,56.5,-43.5</points>
<intersection>35.5 0</intersection>
<intersection>56.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>31.5,-44,35.5,-44</points>
<connection>
<GID>43</GID>
<name>OUT</name></connection>
<intersection>35.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>56.5,-44.5,56.5,-43.5</points>
<connection>
<GID>64</GID>
<name>IN_2</name></connection>
<intersection>-43.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>35.5,-45.5,39.5,-45.5</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-54,35.5,-47.5</points>
<intersection>-54 1</intersection>
<intersection>-50 2</intersection>
<intersection>-47.5 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35.5,-54,56.5,-54</points>
<connection>
<GID>66</GID>
<name>IN_2</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>31.5,-50,35.5,-50</points>
<connection>
<GID>44</GID>
<name>OUT</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>35.5,-47.5,39.5,-47.5</points>
<connection>
<GID>45</GID>
<name>IN_1</name></connection>
<intersection>35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>6.5,-60.5,12.5,-60.5</points>
<connection>
<GID>47</GID>
<name>OUT_0</name></connection>
<connection>
<GID>46</GID>
<name>IN_0</name></connection>
<intersection>9.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>9.5,-64,9.5,-60.5</points>
<intersection>-64 7</intersection>
<intersection>-60.5 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>9.5,-64,26,-64</points>
<intersection>9.5 6</intersection>
<intersection>26 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>26,-66.5,26,-64</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<intersection>-64 7</intersection></vsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>0.5,-69,12.5,-69</points>
<connection>
<GID>48</GID>
<name>OUT_0</name></connection>
<intersection>9.5 6</intersection>
<intersection>12.5 12</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>9.5,-69,9.5,-65</points>
<intersection>-69 1</intersection>
<intersection>-65 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>9.5,-65,24.5,-65</points>
<intersection>9.5 6</intersection>
<intersection>24.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>24.5,-65,24.5,-62.5</points>
<intersection>-65 7</intersection>
<intersection>-62.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>24.5,-62.5,26,-62.5</points>
<connection>
<GID>50</GID>
<name>IN_1</name></connection>
<intersection>24.5 8</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>12.5,-69,12.5,-68.5</points>
<connection>
<GID>49</GID>
<name>IN_0</name></connection>
<intersection>-69 1</intersection></vsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>18.5,-68.5,26,-68.5</points>
<connection>
<GID>51</GID>
<name>IN_1</name></connection>
<connection>
<GID>49</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>18.5,-60.5,26,-60.5</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<connection>
<GID>46</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>32,-61.5,56.5,-61.5</points>
<connection>
<GID>50</GID>
<name>OUT</name></connection>
<intersection>40 4</intersection>
<intersection>56.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>56.5,-62.5,56.5,-61.5</points>
<connection>
<GID>68</GID>
<name>IN_3</name></connection>
<intersection>-61.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>40,-63.5,40,-61.5</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<intersection>-61.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-73,36,-65.5</points>
<intersection>-73 1</intersection>
<intersection>-67.5 2</intersection>
<intersection>-65.5 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,-73,56.5,-73</points>
<connection>
<GID>70</GID>
<name>IN_3</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32,-67.5,36,-67.5</points>
<connection>
<GID>51</GID>
<name>OUT</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>36,-65.5,40,-65.5</points>
<connection>
<GID>52</GID>
<name>IN_1</name></connection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,-76,54,-12.5</points>
<intersection>-76 14</intersection>
<intersection>-67 12</intersection>
<intersection>-56.5 10</intersection>
<intersection>-50 8</intersection>
<intersection>-40.5 6</intersection>
<intersection>-35 4</intersection>
<intersection>-23.5 1</intersection>
<intersection>-12.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54,-23.5,56.5,-23.5</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<intersection>54 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>45.5,-12.5,54,-12.5</points>
<connection>
<GID>31</GID>
<name>OUT</name></connection>
<intersection>54 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>54,-35,56.5,-35</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<intersection>54 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>54,-40.5,56.5,-40.5</points>
<connection>
<GID>64</GID>
<name>IN_0</name></connection>
<intersection>54 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>54,-50,56.5,-50</points>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<intersection>54 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>54,-56.5,56.5,-56.5</points>
<connection>
<GID>68</GID>
<name>IN_0</name></connection>
<intersection>54 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>54,-67,56.5,-67</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>54 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>54,-76,56.5,-76</points>
<connection>
<GID>72</GID>
<name>IN_0</name></connection>
<intersection>54 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,-78,52.5,-29</points>
<intersection>-78 10</intersection>
<intersection>-69 8</intersection>
<intersection>-58.5 6</intersection>
<intersection>-52 4</intersection>
<intersection>-42.5 1</intersection>
<intersection>-29 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52.5,-42.5,56.5,-42.5</points>
<connection>
<GID>64</GID>
<name>IN_1</name></connection>
<intersection>52.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>45.5,-29,52.5,-29</points>
<connection>
<GID>38</GID>
<name>OUT</name></connection>
<intersection>52.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>52.5,-52,56.5,-52</points>
<connection>
<GID>66</GID>
<name>IN_1</name></connection>
<intersection>52.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>52.5,-58.5,56.5,-58.5</points>
<connection>
<GID>68</GID>
<name>IN_1</name></connection>
<intersection>52.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>52.5,-69,56.5,-69</points>
<connection>
<GID>70</GID>
<name>IN_1</name></connection>
<intersection>52.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>52.5,-78,56.5,-78</points>
<connection>
<GID>72</GID>
<name>IN_1</name></connection>
<intersection>52.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51,-80,51,-46.5</points>
<intersection>-80 6</intersection>
<intersection>-71 4</intersection>
<intersection>-60.5 2</intersection>
<intersection>-46.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45.5,-46.5,51,-46.5</points>
<connection>
<GID>45</GID>
<name>OUT</name></connection>
<intersection>51 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>51,-60.5,56.5,-60.5</points>
<connection>
<GID>68</GID>
<name>IN_2</name></connection>
<intersection>51 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>51,-71,56.5,-71</points>
<connection>
<GID>70</GID>
<name>IN_2</name></connection>
<intersection>51 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>51,-80,56.5,-80</points>
<connection>
<GID>72</GID>
<name>IN_2</name></connection>
<intersection>51 0</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,-82,47.5,-64.5</points>
<intersection>-82 1</intersection>
<intersection>-64.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47.5,-82,56.5,-82</points>
<connection>
<GID>72</GID>
<name>IN_3</name></connection>
<intersection>47.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>46,-64.5,47.5,-64.5</points>
<connection>
<GID>52</GID>
<name>OUT</name></connection>
<intersection>47.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75,-79,75,-78.5</points>
<intersection>-79 2</intersection>
<intersection>-78.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>75,-78.5,88,-78.5</points>
<connection>
<GID>84</GID>
<name>N_in0</name></connection>
<intersection>75 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>62.5,-79,75,-79</points>
<connection>
<GID>72</GID>
<name>OUT</name></connection>
<intersection>75 0</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-70,73,-54</points>
<intersection>-70 2</intersection>
<intersection>-54 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73,-54,77,-54</points>
<connection>
<GID>76</GID>
<name>IN_3</name></connection>
<intersection>73 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>62.5,-70,73,-70</points>
<connection>
<GID>70</GID>
<name>OUT</name></connection>
<intersection>73 0</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>62.5,-52,77,-52</points>
<connection>
<GID>66</GID>
<name>OUT</name></connection>
<connection>
<GID>76</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68,-50,68,-36</points>
<intersection>-50 1</intersection>
<intersection>-36 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68,-50,77,-50</points>
<connection>
<GID>76</GID>
<name>IN_1</name></connection>
<intersection>68 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>62.5,-36,68,-36</points>
<connection>
<GID>56</GID>
<name>OUT</name></connection>
<intersection>68 0</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86,-51.5,86,-51</points>
<intersection>-51.5 1</intersection>
<intersection>-51 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>86,-51.5,88,-51.5</points>
<connection>
<GID>82</GID>
<name>N_in0</name></connection>
<intersection>86 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>84,-51,86,-51</points>
<connection>
<GID>76</GID>
<name>OUT</name></connection>
<intersection>86 0</intersection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71.5,-59.5,71.5,-37.5</points>
<intersection>-59.5 2</intersection>
<intersection>-37.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>71.5,-37.5,77,-37.5</points>
<connection>
<GID>74</GID>
<name>IN_3</name></connection>
<intersection>71.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>62.5,-59.5,71.5,-59.5</points>
<connection>
<GID>68</GID>
<name>OUT</name></connection>
<intersection>71.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70.5,-42.5,70.5,-35.5</points>
<intersection>-42.5 2</intersection>
<intersection>-35.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>70.5,-35.5,77,-35.5</points>
<connection>
<GID>74</GID>
<name>IN_2</name></connection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>62.5,-42.5,70.5,-42.5</points>
<connection>
<GID>64</GID>
<name>OUT</name></connection>
<intersection>70.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69.5,-33.5,69.5,-24.5</points>
<intersection>-33.5 1</intersection>
<intersection>-24.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>69.5,-33.5,77,-33.5</points>
<connection>
<GID>74</GID>
<name>IN_1</name></connection>
<intersection>69.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>62.5,-24.5,69.5,-24.5</points>
<connection>
<GID>54</GID>
<name>OUT</name></connection>
<intersection>69.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86,-36,86,-34.5</points>
<intersection>-36 1</intersection>
<intersection>-34.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>86,-36,88,-36</points>
<connection>
<GID>78</GID>
<name>N_in0</name></connection>
<intersection>86 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>84,-34.5,86,-34.5</points>
<connection>
<GID>74</GID>
<name>OUT</name></connection>
<intersection>86 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,62.4,-69.3</PageViewport></page 1>
<page 2>
<PageViewport>0,0,62.4,-69.3</PageViewport></page 2>
<page 3>
<PageViewport>0,0,62.4,-69.3</PageViewport></page 3>
<page 4>
<PageViewport>0,0,62.4,-69.3</PageViewport></page 4>
<page 5>
<PageViewport>0,0,62.4,-69.3</PageViewport></page 5>
<page 6>
<PageViewport>0,0,62.4,-69.3</PageViewport></page 6>
<page 7>
<PageViewport>0,0,62.4,-69.3</PageViewport></page 7>
<page 8>
<PageViewport>0,0,62.4,-69.3</PageViewport></page 8>
<page 9>
<PageViewport>0,0,62.4,-69.3</PageViewport></page 9></circuit>