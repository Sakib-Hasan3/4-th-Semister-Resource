<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>30.4937,1.09687,108.906,-38.3906</PageViewport>
<gate>
<ID>2</ID>
<type>AA_FULLADDER_1BIT</type>
<position>80.5,-17</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_B_0</ID>4 </input>
<output>
<ID>OUT_0</ID>13 </output>
<input>
<ID>carry_in</ID>18 </input>
<output>
<ID>carry_out</ID>1 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3</ID>
<type>AA_FULLADDER_1BIT</type>
<position>71,-17</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_B_0</ID>8 </input>
<output>
<ID>OUT_0</ID>14 </output>
<input>
<ID>carry_in</ID>1 </input>
<output>
<ID>carry_out</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_FULLADDER_1BIT</type>
<position>61.5,-17</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_B_0</ID>10 </input>
<output>
<ID>OUT_0</ID>15 </output>
<input>
<ID>carry_in</ID>2 </input>
<output>
<ID>carry_out</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5</ID>
<type>AA_FULLADDER_1BIT</type>
<position>52,-17</position>
<input>
<ID>IN_0</ID>11 </input>
<input>
<ID>IN_B_0</ID>12 </input>
<output>
<ID>OUT_0</ID>16 </output>
<input>
<ID>carry_in</ID>3 </input>
<output>
<ID>carry_out</ID>17 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7</ID>
<type>GA_LED</type>
<position>52,-23.5</position>
<input>
<ID>N_in3</ID>16 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>9</ID>
<type>GA_LED</type>
<position>46,-23.5</position>
<input>
<ID>N_in3</ID>17 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>11</ID>
<type>GA_LED</type>
<position>61.5,-23.5</position>
<input>
<ID>N_in3</ID>15 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>13</ID>
<type>GA_LED</type>
<position>71,-23.5</position>
<input>
<ID>N_in3</ID>14 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>15</ID>
<type>GA_LED</type>
<position>80.5,-23.5</position>
<input>
<ID>N_in3</ID>13 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>17</ID>
<type>AA_TOGGLE</type>
<position>83,-7</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>19</ID>
<type>AA_TOGGLE</type>
<position>79,-10.5</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_TOGGLE</type>
<position>73,-7</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>21</ID>
<type>AA_TOGGLE</type>
<position>69,-10.5</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_TOGGLE</type>
<position>64,-7</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>23</ID>
<type>AA_TOGGLE</type>
<position>60,-10.5</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_TOGGLE</type>
<position>54,-7</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>25</ID>
<type>AA_TOGGLE</type>
<position>50,-10.5</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>27</ID>
<type>AA_TOGGLE</type>
<position>92.5,-13.5</position>
<output>
<ID>OUT_0</ID>18 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>29</ID>
<type>AA_LABEL</type>
<position>54,-4</position>
<gparam>LABEL_TEXT A3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>30</ID>
<type>AA_LABEL</type>
<position>50,-8</position>
<gparam>LABEL_TEXT B3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>31</ID>
<type>AA_LABEL</type>
<position>60,-8</position>
<gparam>LABEL_TEXT B2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>32</ID>
<type>AA_LABEL</type>
<position>64,-4</position>
<gparam>LABEL_TEXT A2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>33</ID>
<type>AA_LABEL</type>
<position>73,-4</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>34</ID>
<type>AA_LABEL</type>
<position>83,-4</position>
<gparam>LABEL_TEXT A0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>35</ID>
<type>AA_LABEL</type>
<position>79,-8</position>
<gparam>LABEL_TEXT B0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>36</ID>
<type>AA_LABEL</type>
<position>69,-8</position>
<gparam>LABEL_TEXT B1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>37</ID>
<type>AA_LABEL</type>
<position>92.5,-11</position>
<gparam>LABEL_TEXT C in</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>38</ID>
<type>AA_LABEL</type>
<position>80.5,-25.5</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>39</ID>
<type>AA_LABEL</type>
<position>71,-25.5</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>40</ID>
<type>AA_LABEL</type>
<position>61.5,-25.5</position>
<gparam>LABEL_TEXT S2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>41</ID>
<type>AA_LABEL</type>
<position>52,-25.5</position>
<gparam>LABEL_TEXT S3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>42</ID>
<type>AA_LABEL</type>
<position>46,-25.5</position>
<gparam>LABEL_TEXT C4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75,-17,76.5,-17</points>
<connection>
<GID>3</GID>
<name>carry_in</name></connection>
<connection>
<GID>2</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>65.5,-17,67,-17</points>
<connection>
<GID>4</GID>
<name>carry_in</name></connection>
<connection>
<GID>3</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>56,-17,57.5,-17</points>
<connection>
<GID>5</GID>
<name>carry_in</name></connection>
<connection>
<GID>4</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79.5,-14,79.5,-13</points>
<connection>
<GID>2</GID>
<name>IN_B_0</name></connection>
<intersection>-13 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>79,-13,79,-12.5</points>
<connection>
<GID>19</GID>
<name>OUT_0</name></connection>
<intersection>-13 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>79,-13,79.5,-13</points>
<intersection>79 1</intersection>
<intersection>79.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81.5,-14,81.5,-11.5</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>-11.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>83,-11.5,83,-9</points>
<connection>
<GID>17</GID>
<name>OUT_0</name></connection>
<intersection>-11.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>81.5,-11.5,83,-11.5</points>
<intersection>81.5 0</intersection>
<intersection>83 1</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72,-14,72,-11.5</points>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<intersection>-11.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>73,-11.5,73,-9</points>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<intersection>-11.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>72,-11.5,73,-11.5</points>
<intersection>72 0</intersection>
<intersection>73 1</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70,-14,70,-13</points>
<connection>
<GID>3</GID>
<name>IN_B_0</name></connection>
<intersection>-13 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>69,-13,69,-12.5</points>
<connection>
<GID>21</GID>
<name>OUT_0</name></connection>
<intersection>-13 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>69,-13,70,-13</points>
<intersection>69 1</intersection>
<intersection>70 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62.5,-14,62.5,-11.5</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>-11.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>64,-11.5,64,-9</points>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection>
<intersection>-11.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>62.5,-11.5,64,-11.5</points>
<intersection>62.5 0</intersection>
<intersection>64 1</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,-14,60.5,-13</points>
<connection>
<GID>4</GID>
<name>IN_B_0</name></connection>
<intersection>-13 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>60,-13,60,-12.5</points>
<connection>
<GID>23</GID>
<name>OUT_0</name></connection>
<intersection>-13 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>60,-13,60.5,-13</points>
<intersection>60 1</intersection>
<intersection>60.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,-14,53,-11.5</points>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<intersection>-11.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>54,-11.5,54,-9</points>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection>
<intersection>-11.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>53,-11.5,54,-11.5</points>
<intersection>53 0</intersection>
<intersection>54 1</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51,-14,51,-13</points>
<connection>
<GID>5</GID>
<name>IN_B_0</name></connection>
<intersection>-13 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>50,-13,50,-12.5</points>
<connection>
<GID>25</GID>
<name>OUT_0</name></connection>
<intersection>-13 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>50,-13,51,-13</points>
<intersection>50 1</intersection>
<intersection>51 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80.5,-22.5,80.5,-20</points>
<connection>
<GID>15</GID>
<name>N_in3</name></connection>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71,-22.5,71,-20</points>
<connection>
<GID>13</GID>
<name>N_in3</name></connection>
<connection>
<GID>3</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61.5,-22.5,61.5,-20</points>
<connection>
<GID>11</GID>
<name>N_in3</name></connection>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,-22.5,52,-20</points>
<connection>
<GID>7</GID>
<name>N_in3</name></connection>
<connection>
<GID>5</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46,-22.5,46,-17</points>
<connection>
<GID>9</GID>
<name>N_in3</name></connection>
<intersection>-17 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46,-17,48,-17</points>
<connection>
<GID>5</GID>
<name>carry_out</name></connection>
<intersection>46 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>84.5,-13.5,90.5,-13.5</points>
<connection>
<GID>27</GID>
<name>OUT_0</name></connection>
<intersection>84.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>84.5,-17,84.5,-13.5</points>
<connection>
<GID>2</GID>
<name>carry_in</name></connection>
<intersection>-13.5 1</intersection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 1>
<page 2>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 2>
<page 3>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 3>
<page 4>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 4>
<page 5>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 5>
<page 6>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 6>
<page 7>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 7>
<page 8>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 8>
<page 9>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 9></circuit>