<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>0,0,139.4,-70.2</PageViewport>
<gate>
<ID>2</ID>
<type>AA_TOGGLE</type>
<position>11,-5.5</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>11,-8.5</position>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>5</ID>
<type>AA_TOGGLE</type>
<position>11,-11.5</position>
<output>
<ID>OUT_0</ID>23 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>11,-14.5</position>
<output>
<ID>OUT_0</ID>24 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>7</ID>
<type>AA_TOGGLE</type>
<position>11,-18</position>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_TOGGLE</type>
<position>11,-21</position>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>9</ID>
<type>AA_TOGGLE</type>
<position>11,-24</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_TOGGLE</type>
<position>11,-27</position>
<output>
<ID>OUT_0</ID>18 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>11</ID>
<type>AA_TOGGLE</type>
<position>11,-30</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_TOGGLE</type>
<position>11,-33</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>13</ID>
<type>AA_TOGGLE</type>
<position>11,-36</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_TOGGLE</type>
<position>11,-39</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>15</ID>
<type>AA_TOGGLE</type>
<position>11,-42.5</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_TOGGLE</type>
<position>11,-45.5</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>17</ID>
<type>AA_TOGGLE</type>
<position>11,-48.5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_TOGGLE</type>
<position>11,-51.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>20</ID>
<type>DE_OR8</type>
<position>81,-14</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>7 </input>
<input>
<ID>IN_2</ID>6 </input>
<input>
<ID>IN_3</ID>5 </input>
<input>
<ID>IN_4</ID>1 </input>
<input>
<ID>IN_5</ID>2 </input>
<input>
<ID>IN_6</ID>3 </input>
<input>
<ID>IN_7</ID>4 </input>
<output>
<ID>OUT</ID>26 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>24</ID>
<type>DE_OR8</type>
<position>81,-24</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>16 </input>
<input>
<ID>IN_2</ID>17 </input>
<input>
<ID>IN_3</ID>18 </input>
<input>
<ID>IN_4</ID>1 </input>
<input>
<ID>IN_5</ID>2 </input>
<input>
<ID>IN_6</ID>3 </input>
<input>
<ID>IN_7</ID>4 </input>
<output>
<ID>OUT</ID>27 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>25</ID>
<type>DE_OR8</type>
<position>81,-34.5</position>
<input>
<ID>IN_0</ID>23 </input>
<input>
<ID>IN_1</ID>24 </input>
<input>
<ID>IN_2</ID>17 </input>
<input>
<ID>IN_3</ID>18 </input>
<input>
<ID>IN_4</ID>1 </input>
<input>
<ID>IN_5</ID>2 </input>
<input>
<ID>IN_6</ID>5 </input>
<input>
<ID>IN_7</ID>6 </input>
<output>
<ID>OUT</ID>28 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>26</ID>
<type>DE_OR8</type>
<position>81,-44.5</position>
<input>
<ID>IN_0</ID>25 </input>
<input>
<ID>IN_1</ID>24 </input>
<input>
<ID>IN_2</ID>16 </input>
<input>
<ID>IN_3</ID>18 </input>
<input>
<ID>IN_4</ID>1 </input>
<input>
<ID>IN_5</ID>3 </input>
<input>
<ID>IN_6</ID>5 </input>
<input>
<ID>IN_7</ID>7 </input>
<output>
<ID>OUT</ID>29 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>28</ID>
<type>GA_LED</type>
<position>90,-14</position>
<input>
<ID>N_in0</ID>26 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>29</ID>
<type>GA_LED</type>
<position>90,-24.5</position>
<input>
<ID>N_in0</ID>27 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>30</ID>
<type>GA_LED</type>
<position>90,-35</position>
<input>
<ID>N_in0</ID>28 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>31</ID>
<type>GA_LED</type>
<position>90,-45.5</position>
<input>
<ID>N_in0</ID>29 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42.5,-51,42.5,-17.5</points>
<intersection>-51 2</intersection>
<intersection>-17.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>42.5,-17.5,78,-17.5</points>
<connection>
<GID>20</GID>
<name>IN_4</name></connection>
<intersection>42.5 0</intersection>
<intersection>73.5 5</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13.5,-51,42.5,-51</points>
<intersection>13.5 3</intersection>
<intersection>42.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>13.5,-51.5,13.5,-51</points>
<intersection>-51.5 4</intersection>
<intersection>-51 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>13,-51.5,13.5,-51.5</points>
<connection>
<GID>18</GID>
<name>OUT_0</name></connection>
<intersection>13.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>73.5,-27.5,73.5,-17.5</points>
<intersection>-27.5 6</intersection>
<intersection>-17.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>72,-27.5,78,-27.5</points>
<connection>
<GID>24</GID>
<name>IN_4</name></connection>
<intersection>72 7</intersection>
<intersection>73.5 5</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>72,-38,72,-27.5</points>
<intersection>-38 8</intersection>
<intersection>-27.5 6</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>72,-38,78,-38</points>
<connection>
<GID>25</GID>
<name>IN_4</name></connection>
<intersection>72 7</intersection>
<intersection>74.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>74.5,-48,74.5,-38</points>
<intersection>-48 10</intersection>
<intersection>-38 8</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>74.5,-48,78,-48</points>
<connection>
<GID>26</GID>
<name>IN_4</name></connection>
<intersection>74.5 9</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,-48.5,40.5,-16.5</points>
<intersection>-48.5 2</intersection>
<intersection>-16.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40.5,-16.5,78,-16.5</points>
<connection>
<GID>20</GID>
<name>IN_5</name></connection>
<intersection>40.5 0</intersection>
<intersection>74.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13,-48.5,40.5,-48.5</points>
<connection>
<GID>17</GID>
<name>OUT_0</name></connection>
<intersection>40.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>74.5,-26.5,74.5,-16.5</points>
<intersection>-26.5 4</intersection>
<intersection>-16.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>74.5,-26.5,78,-26.5</points>
<connection>
<GID>24</GID>
<name>IN_5</name></connection>
<intersection>74.5 3</intersection>
<intersection>75.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>75.5,-37,75.5,-26.5</points>
<intersection>-37 6</intersection>
<intersection>-26.5 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>75.5,-37,78,-37</points>
<connection>
<GID>25</GID>
<name>IN_5</name></connection>
<intersection>75.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-52,39,-15.5</points>
<intersection>-52 2</intersection>
<intersection>-15.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39,-15.5,78,-15.5</points>
<connection>
<GID>20</GID>
<name>IN_6</name></connection>
<intersection>39 0</intersection>
<intersection>76 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34.5,-52,39,-52</points>
<intersection>34.5 5</intersection>
<intersection>39 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>34.5,-52,34.5,-45.5</points>
<intersection>-52 2</intersection>
<intersection>-45.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>13,-45.5,34.5,-45.5</points>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection>
<intersection>34.5 5</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>76,-25.5,76,-15.5</points>
<intersection>-25.5 8</intersection>
<intersection>-15.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>68,-25.5,78,-25.5</points>
<connection>
<GID>24</GID>
<name>IN_6</name></connection>
<intersection>68 9</intersection>
<intersection>76 7</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>68,-47,68,-25.5</points>
<intersection>-47 10</intersection>
<intersection>-25.5 8</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>68,-47,78,-47</points>
<connection>
<GID>26</GID>
<name>IN_5</name></connection>
<intersection>68 9</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,-42.5,38,-14.5</points>
<intersection>-42.5 2</intersection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38,-14.5,78,-14.5</points>
<connection>
<GID>20</GID>
<name>IN_7</name></connection>
<intersection>38 0</intersection>
<intersection>77 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13,-42.5,38,-42.5</points>
<connection>
<GID>15</GID>
<name>OUT_0</name></connection>
<intersection>38 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>77,-24.5,77,-14.5</points>
<intersection>-24.5 4</intersection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>77,-24.5,78,-24.5</points>
<connection>
<GID>24</GID>
<name>IN_7</name></connection>
<intersection>77 3</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35.5,-13.5,78,-13.5</points>
<connection>
<GID>20</GID>
<name>IN_3</name></connection>
<intersection>35.5 3</intersection>
<intersection>69.5 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>35.5,-39,35.5,-13.5</points>
<intersection>-39 4</intersection>
<intersection>-13.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>13,-39,35.5,-39</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>35.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>69.5,-36,69.5,-13.5</points>
<intersection>-36 6</intersection>
<intersection>-13.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>63.5,-36,78,-36</points>
<connection>
<GID>25</GID>
<name>IN_6</name></connection>
<intersection>63.5 7</intersection>
<intersection>69.5 5</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>63.5,-46,63.5,-36</points>
<intersection>-46 8</intersection>
<intersection>-36 6</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>63.5,-46,78,-46</points>
<connection>
<GID>26</GID>
<name>IN_6</name></connection>
<intersection>63.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37.5,-36,37.5,-12.5</points>
<intersection>-36 2</intersection>
<intersection>-12.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37.5,-12.5,78,-12.5</points>
<connection>
<GID>20</GID>
<name>IN_2</name></connection>
<intersection>37.5 0</intersection>
<intersection>66 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13,-36,37.5,-36</points>
<connection>
<GID>13</GID>
<name>OUT_0</name></connection>
<intersection>37.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>66,-35,66,-12.5</points>
<intersection>-35 4</intersection>
<intersection>-12.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>66,-35,78,-35</points>
<connection>
<GID>25</GID>
<name>IN_7</name></connection>
<intersection>66 3</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36.5,-33,36.5,-11.5</points>
<intersection>-33 2</intersection>
<intersection>-11.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36.5,-11.5,78,-11.5</points>
<connection>
<GID>20</GID>
<name>IN_1</name></connection>
<intersection>36.5 0</intersection>
<intersection>70.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13,-33,36.5,-33</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<intersection>36.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>70.5,-45,70.5,-11.5</points>
<intersection>-45 4</intersection>
<intersection>-11.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>70.5,-45,78,-45</points>
<connection>
<GID>26</GID>
<name>IN_7</name></connection>
<intersection>70.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-30,39,-10.5</points>
<intersection>-30 2</intersection>
<intersection>-10.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39,-10.5,78,-10.5</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13,-30,39,-30</points>
<connection>
<GID>11</GID>
<name>OUT_0</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45.5,-20.5,45.5,-18</points>
<intersection>-20.5 1</intersection>
<intersection>-18 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45.5,-20.5,78,-20.5</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>45.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13,-18,45.5,-18</points>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection>
<intersection>45.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45.5,-21.5,45.5,-21</points>
<intersection>-21.5 1</intersection>
<intersection>-21 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45.5,-21.5,78,-21.5</points>
<connection>
<GID>24</GID>
<name>IN_1</name></connection>
<intersection>45.5 0</intersection>
<intersection>70.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13,-21,45.5,-21</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>45.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>70.5,-43,70.5,-21.5</points>
<intersection>-43 4</intersection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>70.5,-43,78,-43</points>
<connection>
<GID>26</GID>
<name>IN_2</name></connection>
<intersection>70.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45.5,-24,45.5,-22.5</points>
<intersection>-24 2</intersection>
<intersection>-22.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45.5,-22.5,78,-22.5</points>
<connection>
<GID>24</GID>
<name>IN_2</name></connection>
<intersection>45.5 0</intersection>
<intersection>74.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13,-24,45.5,-24</points>
<connection>
<GID>9</GID>
<name>OUT_0</name></connection>
<intersection>45.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>74.5,-33,74.5,-22.5</points>
<intersection>-33 4</intersection>
<intersection>-22.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>74.5,-33,78,-33</points>
<connection>
<GID>25</GID>
<name>IN_2</name></connection>
<intersection>74.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48.5,-27,48.5,-23.5</points>
<intersection>-27 2</intersection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>48.5,-23.5,78,-23.5</points>
<connection>
<GID>24</GID>
<name>IN_3</name></connection>
<intersection>48.5 0</intersection>
<intersection>77 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13,-27,48.5,-27</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>48.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>77,-34,77,-23.5</points>
<intersection>-34 4</intersection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>73.5,-34,78,-34</points>
<connection>
<GID>25</GID>
<name>IN_3</name></connection>
<intersection>73.5 5</intersection>
<intersection>77 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>73.5,-44,73.5,-34</points>
<intersection>-44 6</intersection>
<intersection>-34 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>73.5,-44,78,-44</points>
<connection>
<GID>26</GID>
<name>IN_3</name></connection>
<intersection>73.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,-31,47.5,-11.5</points>
<intersection>-31 1</intersection>
<intersection>-11.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47.5,-31,78,-31</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>47.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13,-11.5,47.5,-11.5</points>
<connection>
<GID>5</GID>
<name>OUT_0</name></connection>
<intersection>47.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45.5,-32,45.5,-14.5</points>
<intersection>-32 1</intersection>
<intersection>-14.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45.5,-32,78,-32</points>
<connection>
<GID>25</GID>
<name>IN_1</name></connection>
<intersection>45.5 0</intersection>
<intersection>72.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13,-14.5,45.5,-14.5</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>45.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>72.5,-42,72.5,-32</points>
<intersection>-42 4</intersection>
<intersection>-32 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>72.5,-42,78,-42</points>
<connection>
<GID>26</GID>
<name>IN_1</name></connection>
<intersection>72.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45.5,-41,45.5,-8.5</points>
<intersection>-41 2</intersection>
<intersection>-8.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>13,-8.5,45.5,-8.5</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>45.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>45.5,-41,78,-41</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>45.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>85,-14,89,-14</points>
<connection>
<GID>28</GID>
<name>N_in0</name></connection>
<connection>
<GID>20</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87,-24.5,87,-24</points>
<intersection>-24.5 1</intersection>
<intersection>-24 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>87,-24.5,89,-24.5</points>
<connection>
<GID>29</GID>
<name>N_in0</name></connection>
<intersection>87 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>85,-24,87,-24</points>
<connection>
<GID>24</GID>
<name>OUT</name></connection>
<intersection>87 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87,-35,87,-34.5</points>
<intersection>-35 1</intersection>
<intersection>-34.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>87,-35,89,-35</points>
<connection>
<GID>30</GID>
<name>N_in0</name></connection>
<intersection>87 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>85,-34.5,87,-34.5</points>
<connection>
<GID>25</GID>
<name>OUT</name></connection>
<intersection>87 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87,-45.5,87,-44.5</points>
<intersection>-45.5 1</intersection>
<intersection>-44.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>87,-45.5,89,-45.5</points>
<connection>
<GID>31</GID>
<name>N_in0</name></connection>
<intersection>87 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>85,-44.5,87,-44.5</points>
<connection>
<GID>26</GID>
<name>OUT</name></connection>
<intersection>87 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 1>
<page 2>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 2>
<page 3>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 3>
<page 4>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 4>
<page 5>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 5>
<page 6>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 6>
<page 7>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 7>
<page 8>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 8>
<page 9>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 9></circuit>