<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>0,0,139.4,-70.2</PageViewport>
<gate>
<ID>2</ID>
<type>AA_FULLADDER_1BIT</type>
<position>29,-15</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_B_0</ID>11 </input>
<output>
<ID>OUT_0</ID>12 </output>
<input>
<ID>carry_in</ID>3 </input>
<output>
<ID>carry_out</ID>16 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_FULLADDER_1BIT</type>
<position>38,-15</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_B_0</ID>9 </input>
<output>
<ID>OUT_0</ID>13 </output>
<input>
<ID>carry_in</ID>1 </input>
<output>
<ID>carry_out</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5</ID>
<type>AA_FULLADDER_1BIT</type>
<position>46.5,-15</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_B_0</ID>7 </input>
<output>
<ID>OUT_0</ID>14 </output>
<input>
<ID>carry_in</ID>2 </input>
<output>
<ID>carry_out</ID>1 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_FULLADDER_1BIT</type>
<position>55.5,-15</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_B_0</ID>5 </input>
<output>
<ID>OUT_0</ID>15 </output>
<output>
<ID>carry_out</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_TOGGLE</type>
<position>45,-3.5</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_TOGGLE</type>
<position>47.5,-3.5</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>11</ID>
<type>AA_TOGGLE</type>
<position>55,-4</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_TOGGLE</type>
<position>57.5,-4</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>13</ID>
<type>AA_TOGGLE</type>
<position>36.5,-4</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_TOGGLE</type>
<position>39,-4</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>15</ID>
<type>AA_TOGGLE</type>
<position>28,-4</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_TOGGLE</type>
<position>30.5,-4</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>18</ID>
<type>GA_LED</type>
<position>28,-25</position>
<input>
<ID>N_in3</ID>12 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>19</ID>
<type>GA_LED</type>
<position>37.5,-26</position>
<input>
<ID>N_in3</ID>13 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>GA_LED</type>
<position>46.5,-26</position>
<input>
<ID>N_in3</ID>14 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>21</ID>
<type>GA_LED</type>
<position>55.5,-26.5</position>
<input>
<ID>N_in3</ID>15 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>23</ID>
<type>GA_LED</type>
<position>19.5,-15.5</position>
<input>
<ID>N_in1</ID>16 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>42,-15,42.5,-15</points>
<connection>
<GID>4</GID>
<name>carry_in</name></connection>
<connection>
<GID>5</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50.5,-15,51.5,-15</points>
<connection>
<GID>5</GID>
<name>carry_in</name></connection>
<connection>
<GID>6</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33,-15,34,-15</points>
<connection>
<GID>4</GID>
<name>carry_out</name></connection>
<connection>
<GID>2</GID>
<name>carry_in</name></connection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,-12,56.5,-9</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>-9 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>57.5,-9,57.5,-6</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<intersection>-9 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>56.5,-9,57.5,-9</points>
<intersection>56.5 0</intersection>
<intersection>57.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-12,54.5,-9</points>
<connection>
<GID>6</GID>
<name>IN_B_0</name></connection>
<intersection>-9 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>55,-9,55,-6</points>
<connection>
<GID>11</GID>
<name>OUT_0</name></connection>
<intersection>-9 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>54.5,-9,55,-9</points>
<intersection>54.5 0</intersection>
<intersection>55 1</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,-12,47.5,-5.5</points>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45.5,-12,45.5,-8.5</points>
<connection>
<GID>5</GID>
<name>IN_B_0</name></connection>
<intersection>-8.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>45,-8.5,45,-5.5</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>-8.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>45,-8.5,45.5,-8.5</points>
<intersection>45 1</intersection>
<intersection>45.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-12,39,-6</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-12,37,-9</points>
<connection>
<GID>4</GID>
<name>IN_B_0</name></connection>
<intersection>-9 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>36.5,-9,36.5,-6</points>
<connection>
<GID>13</GID>
<name>OUT_0</name></connection>
<intersection>-9 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>36.5,-9,37,-9</points>
<intersection>36.5 1</intersection>
<intersection>37 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,-12,30,-9</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>-9 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>30.5,-9,30.5,-6</points>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection>
<intersection>-9 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>30,-9,30.5,-9</points>
<intersection>30 0</intersection>
<intersection>30.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-12,28,-6</points>
<connection>
<GID>2</GID>
<name>IN_B_0</name></connection>
<connection>
<GID>15</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-24,28,-21</points>
<connection>
<GID>18</GID>
<name>N_in3</name></connection>
<intersection>-21 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>29,-21,29,-18</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>-21 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>28,-21,29,-21</points>
<intersection>28 0</intersection>
<intersection>29 1</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37.5,-25,37.5,-21.5</points>
<connection>
<GID>19</GID>
<name>N_in3</name></connection>
<intersection>-21.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>38,-21.5,38,-18</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>-21.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>37.5,-21.5,38,-21.5</points>
<intersection>37.5 0</intersection>
<intersection>38 1</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46.5,-25,46.5,-18</points>
<connection>
<GID>20</GID>
<name>N_in3</name></connection>
<connection>
<GID>5</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55.5,-25.5,55.5,-18</points>
<connection>
<GID>21</GID>
<name>N_in3</name></connection>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-15.5,22.5,-15</points>
<intersection>-15.5 2</intersection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22.5,-15,25,-15</points>
<connection>
<GID>2</GID>
<name>carry_out</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>20.5,-15.5,22.5,-15.5</points>
<connection>
<GID>23</GID>
<name>N_in1</name></connection>
<intersection>22.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 1>
<page 2>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 2>
<page 3>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 3>
<page 4>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 4>
<page 5>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 5>
<page 6>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 6>
<page 7>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 7>
<page 8>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 8>
<page 9>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 9></circuit>