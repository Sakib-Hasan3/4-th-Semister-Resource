<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>9.425,9.225,113.975,-43.425</PageViewport>
<gate>
<ID>2</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>44.5,-19</position>
<output>
<ID>A_equal_B</ID>10 </output>
<output>
<ID>A_greater_B</ID>9 </output>
<output>
<ID>A_less_B</ID>11 </output>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>6 </input>
<input>
<ID>IN_2</ID>7 </input>
<input>
<ID>IN_3</ID>8 </input>
<input>
<ID>IN_B_0</ID>4 </input>
<input>
<ID>IN_B_1</ID>3 </input>
<input>
<ID>IN_B_2</ID>2 </input>
<input>
<ID>IN_B_3</ID>1 </input>
<input>
<ID>in_A_equal_B</ID>15 </input>
<input>
<ID>in_A_greater_B</ID>14 </input>
<input>
<ID>in_A_less_B</ID>16 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>49,-7</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>5</ID>
<type>AA_TOGGLE</type>
<position>46.5,-7</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>53.5,-7</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>7</ID>
<type>AA_TOGGLE</type>
<position>51,-7</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_TOGGLE</type>
<position>38.5,-6.5</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>11</ID>
<type>AA_TOGGLE</type>
<position>36,-6.5</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_TOGGLE</type>
<position>43.5,-6.5</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>13</ID>
<type>AA_TOGGLE</type>
<position>40.5,-6.5</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>15</ID>
<type>GA_LED</type>
<position>31.5,-17</position>
<input>
<ID>N_in1</ID>9 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>17</ID>
<type>GA_LED</type>
<position>31.5,-20</position>
<input>
<ID>N_in1</ID>10 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>19</ID>
<type>GA_LED</type>
<position>31.5,-23.5</position>
<input>
<ID>N_in1</ID>11 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>21</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>68.5,-18.5</position>
<output>
<ID>A_equal_B</ID>15 </output>
<output>
<ID>A_greater_B</ID>14 </output>
<output>
<ID>A_less_B</ID>16 </output>
<input>
<ID>IN_0</ID>24 </input>
<input>
<ID>IN_1</ID>23 </input>
<input>
<ID>IN_2</ID>22 </input>
<input>
<ID>IN_3</ID>21 </input>
<input>
<ID>IN_B_0</ID>20 </input>
<input>
<ID>IN_B_1</ID>19 </input>
<input>
<ID>IN_B_2</ID>18 </input>
<input>
<ID>IN_B_3</ID>17 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_TOGGLE</type>
<position>73,-7.5</position>
<output>
<ID>OUT_0</ID>18 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>23</ID>
<type>AA_TOGGLE</type>
<position>70.5,-7.5</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_TOGGLE</type>
<position>77.5,-7.5</position>
<output>
<ID>OUT_0</ID>20 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>25</ID>
<type>AA_TOGGLE</type>
<position>75,-7.5</position>
<output>
<ID>OUT_0</ID>19 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_TOGGLE</type>
<position>62.5,-7</position>
<output>
<ID>OUT_0</ID>22 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>27</ID>
<type>AA_TOGGLE</type>
<position>60,-7</position>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_TOGGLE</type>
<position>67,-7</position>
<output>
<ID>OUT_0</ID>24 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>29</ID>
<type>AA_TOGGLE</type>
<position>64.5,-7</position>
<output>
<ID>OUT_0</ID>23 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46.5,-15,46.5,-9</points>
<connection>
<GID>2</GID>
<name>IN_B_3</name></connection>
<connection>
<GID>5</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,-15,47.5,-12</points>
<connection>
<GID>2</GID>
<name>IN_B_2</name></connection>
<intersection>-12 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>49,-12,49,-9</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>-12 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>47.5,-12,49,-12</points>
<intersection>47.5 0</intersection>
<intersection>49 1</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48.5,-15,48.5,-13</points>
<connection>
<GID>2</GID>
<name>IN_B_1</name></connection>
<intersection>-13 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>51,-13,51,-9</points>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection>
<intersection>-13 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-13,51,-13</points>
<intersection>48.5 0</intersection>
<intersection>51 1</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-15,49.5,-14</points>
<connection>
<GID>2</GID>
<name>IN_B_0</name></connection>
<intersection>-14 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>53.5,-14,53.5,-9</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>-14 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>49.5,-14,53.5,-14</points>
<intersection>49.5 0</intersection>
<intersection>53.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42.5,-15,42.5,-11.5</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>-11.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>43.5,-11.5,43.5,-8.5</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<intersection>-11.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>42.5,-11.5,43.5,-11.5</points>
<intersection>42.5 0</intersection>
<intersection>43.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41.5,-15,41.5,-11.5</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>-11.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>40.5,-11.5,40.5,-8.5</points>
<connection>
<GID>13</GID>
<name>OUT_0</name></connection>
<intersection>-11.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>40.5,-11.5,41.5,-11.5</points>
<intersection>40.5 1</intersection>
<intersection>41.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,-15,40.5,-12</points>
<connection>
<GID>2</GID>
<name>IN_2</name></connection>
<intersection>-12 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>38.5,-12,38.5,-8.5</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>-12 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>38.5,-12,40.5,-12</points>
<intersection>38.5 1</intersection>
<intersection>40.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39.5,-15,39.5,-12.5</points>
<connection>
<GID>2</GID>
<name>IN_3</name></connection>
<intersection>-12.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>36,-12.5,36,-8.5</points>
<connection>
<GID>11</GID>
<name>OUT_0</name></connection>
<intersection>-12.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>36,-12.5,39.5,-12.5</points>
<intersection>36 1</intersection>
<intersection>39.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>32.5,-17,36.5,-17</points>
<connection>
<GID>2</GID>
<name>A_greater_B</name></connection>
<connection>
<GID>15</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,-20,34.5,-19</points>
<intersection>-20 2</intersection>
<intersection>-19 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34.5,-19,36.5,-19</points>
<connection>
<GID>2</GID>
<name>A_equal_B</name></connection>
<intersection>34.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32.5,-20,34.5,-20</points>
<connection>
<GID>17</GID>
<name>N_in1</name></connection>
<intersection>34.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,-23.5,34.5,-21</points>
<intersection>-23.5 2</intersection>
<intersection>-21 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34.5,-21,36.5,-21</points>
<connection>
<GID>2</GID>
<name>A_less_B</name></connection>
<intersection>34.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32.5,-23.5,34.5,-23.5</points>
<connection>
<GID>19</GID>
<name>N_in1</name></connection>
<intersection>34.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,-17,56.5,-16.5</points>
<intersection>-17 4</intersection>
<intersection>-16.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>56.5,-16.5,60.5,-16.5</points>
<connection>
<GID>21</GID>
<name>A_greater_B</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>52.5,-17,56.5,-17</points>
<connection>
<GID>2</GID>
<name>in_A_greater_B</name></connection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,-19,56.5,-18.5</points>
<intersection>-19 4</intersection>
<intersection>-18.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>56.5,-18.5,60.5,-18.5</points>
<connection>
<GID>21</GID>
<name>A_equal_B</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>52.5,-19,56.5,-19</points>
<connection>
<GID>2</GID>
<name>in_A_equal_B</name></connection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,-21,56.5,-20.5</points>
<intersection>-21 4</intersection>
<intersection>-20.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>56.5,-20.5,60.5,-20.5</points>
<connection>
<GID>21</GID>
<name>A_less_B</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>52.5,-21,56.5,-21</points>
<connection>
<GID>2</GID>
<name>in_A_less_B</name></connection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70.5,-14.5,70.5,-9.5</points>
<connection>
<GID>21</GID>
<name>IN_B_3</name></connection>
<connection>
<GID>23</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71.5,-14.5,71.5,-12</points>
<connection>
<GID>21</GID>
<name>IN_B_2</name></connection>
<intersection>-12 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>73,-12,73,-9.5</points>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection>
<intersection>-12 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>71.5,-12,73,-12</points>
<intersection>71.5 0</intersection>
<intersection>73 1</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72.5,-14.5,72.5,-12.5</points>
<connection>
<GID>21</GID>
<name>IN_B_1</name></connection>
<intersection>-12.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>75,-12.5,75,-9.5</points>
<connection>
<GID>25</GID>
<name>OUT_0</name></connection>
<intersection>-12.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>72.5,-12.5,75,-12.5</points>
<intersection>72.5 0</intersection>
<intersection>75 1</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73.5,-14.5,73.5,-13.5</points>
<connection>
<GID>21</GID>
<name>IN_B_0</name></connection>
<intersection>-13.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>77.5,-13.5,77.5,-9.5</points>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection>
<intersection>-13.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>73.5,-13.5,77.5,-13.5</points>
<intersection>73.5 0</intersection>
<intersection>77.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63.5,-14.5,63.5,-12</points>
<connection>
<GID>21</GID>
<name>IN_3</name></connection>
<intersection>-12 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>60,-12,60,-9</points>
<connection>
<GID>27</GID>
<name>OUT_0</name></connection>
<intersection>-12 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>60,-12,63.5,-12</points>
<intersection>60 1</intersection>
<intersection>63.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64.5,-14.5,64.5,-11.5</points>
<connection>
<GID>21</GID>
<name>IN_2</name></connection>
<intersection>-11.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>62.5,-11.5,62.5,-9</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<intersection>-11.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>62.5,-11.5,64.5,-11.5</points>
<intersection>62.5 1</intersection>
<intersection>64.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65.5,-14.5,65.5,-11.5</points>
<connection>
<GID>21</GID>
<name>IN_1</name></connection>
<intersection>-11.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>65,-11.5,65,-9</points>
<intersection>-11.5 2</intersection>
<intersection>-9 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>65,-11.5,65.5,-11.5</points>
<intersection>65 1</intersection>
<intersection>65.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>64.5,-9,65,-9</points>
<connection>
<GID>29</GID>
<name>OUT_0</name></connection>
<intersection>65 1</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67,-11.5,67,-9</points>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection>
<intersection>-11.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>66.5,-14.5,66.5,-11.5</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<intersection>-11.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>66.5,-11.5,67,-11.5</points>
<intersection>66.5 1</intersection>
<intersection>67 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 1>
<page 2>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 2>
<page 3>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 3>
<page 4>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 4>
<page 5>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 5>
<page 6>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 6>
<page 7>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 7>
<page 8>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 8>
<page 9>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 9></circuit>