<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-6.34154,19.5695,159.06,-63.7244</PageViewport>
<gate>
<ID>1</ID>
<type>AE_FULLADDER_4BIT</type>
<position>94.5,-11</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>10 </input>
<input>
<ID>IN_2</ID>11 </input>
<input>
<ID>IN_3</ID>12 </input>
<input>
<ID>IN_B_0</ID>8 </input>
<input>
<ID>IN_B_1</ID>7 </input>
<input>
<ID>IN_B_2</ID>6 </input>
<input>
<ID>IN_B_3</ID>5 </input>
<output>
<ID>OUT_0</ID>4 </output>
<output>
<ID>OUT_1</ID>3 </output>
<output>
<ID>OUT_2</ID>2 </output>
<output>
<ID>OUT_3</ID>1 </output>
<output>
<ID>carry_out</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>2</ID>
<type>AE_FULLADDER_4BIT</type>
<position>91,-41</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>46 </input>
<input>
<ID>IN_2</ID>46 </input>
<input>
<ID>IN_3</ID>17 </input>
<input>
<ID>IN_B_0</ID>4 </input>
<input>
<ID>IN_B_1</ID>3 </input>
<input>
<ID>IN_B_2</ID>2 </input>
<input>
<ID>IN_B_3</ID>1 </input>
<output>
<ID>OUT_0</ID>21 </output>
<output>
<ID>OUT_1</ID>20 </output>
<output>
<ID>OUT_2</ID>19 </output>
<output>
<ID>OUT_3</ID>18 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>3</ID>
<type>AA_TOGGLE</type>
<position>97,9.5</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>99,9.5</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>5</ID>
<type>AA_TOGGLE</type>
<position>101,9.5</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>103,9.5</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>7</ID>
<type>AA_TOGGLE</type>
<position>87.5,9.5</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_TOGGLE</type>
<position>89.5,9.5</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>9</ID>
<type>AA_TOGGLE</type>
<position>91.5,9.5</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_TOGGLE</type>
<position>93.5,9.5</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>11</ID>
<type>AE_OR3</type>
<position>77.5,-16</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>14 </input>
<input>
<ID>IN_2</ID>13 </input>
<output>
<ID>OUT</ID>46 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_AND2</type>
<position>86.5,-17</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>1 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>13</ID>
<type>AA_AND2</type>
<position>86.5,-22</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>1 </input>
<output>
<ID>OUT</ID>15 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>14</ID>
<type>GA_LED</type>
<position>93.5,-49.5</position>
<input>
<ID>N_in3</ID>21 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>15</ID>
<type>GA_LED</type>
<position>91,-49.5</position>
<input>
<ID>N_in3</ID>20 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>16</ID>
<type>GA_LED</type>
<position>88.5,-49.5</position>
<input>
<ID>N_in3</ID>19 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>17</ID>
<type>GA_LED</type>
<position>86,-49.5</position>
<input>
<ID>N_in3</ID>18 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>AE_FULLADDER_4BIT</type>
<position>54,-9.5</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>32 </input>
<input>
<ID>IN_2</ID>33 </input>
<input>
<ID>IN_3</ID>34 </input>
<input>
<ID>IN_B_0</ID>30 </input>
<input>
<ID>IN_B_1</ID>29 </input>
<input>
<ID>IN_B_2</ID>28 </input>
<input>
<ID>IN_B_3</ID>27 </input>
<output>
<ID>OUT_0</ID>26 </output>
<output>
<ID>OUT_1</ID>25 </output>
<output>
<ID>OUT_2</ID>24 </output>
<output>
<ID>OUT_3</ID>23 </output>
<input>
<ID>carry_in</ID>46 </input>
<output>
<ID>carry_out</ID>35 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>21</ID>
<type>AE_FULLADDER_4BIT</type>
<position>50.5,-39.5</position>
<input>
<ID>IN_0</ID>39 </input>
<input>
<ID>IN_1</ID>38 </input>
<input>
<ID>IN_2</ID>38 </input>
<input>
<ID>IN_3</ID>39 </input>
<input>
<ID>IN_B_0</ID>26 </input>
<input>
<ID>IN_B_1</ID>25 </input>
<input>
<ID>IN_B_2</ID>24 </input>
<input>
<ID>IN_B_3</ID>23 </input>
<output>
<ID>OUT_0</ID>43 </output>
<output>
<ID>OUT_1</ID>42 </output>
<output>
<ID>OUT_2</ID>41 </output>
<output>
<ID>OUT_3</ID>40 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_TOGGLE</type>
<position>56.5,11</position>
<output>
<ID>OUT_0</ID>27 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>23</ID>
<type>AA_TOGGLE</type>
<position>58.5,11</position>
<output>
<ID>OUT_0</ID>28 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_TOGGLE</type>
<position>60.5,11</position>
<output>
<ID>OUT_0</ID>29 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>25</ID>
<type>AA_TOGGLE</type>
<position>62.5,11</position>
<output>
<ID>OUT_0</ID>30 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_TOGGLE</type>
<position>47,11</position>
<output>
<ID>OUT_0</ID>34 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>27</ID>
<type>AA_TOGGLE</type>
<position>49,11</position>
<output>
<ID>OUT_0</ID>33 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_TOGGLE</type>
<position>51,11</position>
<output>
<ID>OUT_0</ID>32 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>29</ID>
<type>AA_TOGGLE</type>
<position>53,11</position>
<output>
<ID>OUT_0</ID>31 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>30</ID>
<type>AE_OR3</type>
<position>37,-14.5</position>
<input>
<ID>IN_0</ID>37 </input>
<input>
<ID>IN_1</ID>36 </input>
<input>
<ID>IN_2</ID>35 </input>
<output>
<ID>OUT</ID>38 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>31</ID>
<type>AA_AND2</type>
<position>46,-15.5</position>
<input>
<ID>IN_0</ID>24 </input>
<input>
<ID>IN_1</ID>23 </input>
<output>
<ID>OUT</ID>36 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>32</ID>
<type>AA_AND2</type>
<position>46,-20.5</position>
<input>
<ID>IN_0</ID>25 </input>
<input>
<ID>IN_1</ID>23 </input>
<output>
<ID>OUT</ID>37 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>33</ID>
<type>GA_LED</type>
<position>53,-48</position>
<input>
<ID>N_in3</ID>43 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>GA_LED</type>
<position>50.5,-48</position>
<input>
<ID>N_in3</ID>42 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>35</ID>
<type>GA_LED</type>
<position>48,-48</position>
<input>
<ID>N_in3</ID>41 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>36</ID>
<type>GA_LED</type>
<position>45.5,-48</position>
<input>
<ID>N_in3</ID>40 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>37</ID>
<type>GA_LED</type>
<position>39.5,-47.5</position>
<input>
<ID>N_in3</ID>38 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93,-37,93,-15</points>
<connection>
<GID>2</GID>
<name>IN_B_3</name></connection>
<connection>
<GID>1</GID>
<name>OUT_3</name></connection>
<intersection>-21 7</intersection>
<intersection>-16 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>89.5,-16,93,-16</points>
<connection>
<GID>12</GID>
<name>IN_1</name></connection>
<intersection>93 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>89.5,-21,93,-21</points>
<connection>
<GID>13</GID>
<name>IN_1</name></connection>
<intersection>93 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>94,-37,94,-15</points>
<connection>
<GID>2</GID>
<name>IN_B_2</name></connection>
<connection>
<GID>1</GID>
<name>OUT_2</name></connection>
<intersection>-18 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>89.5,-18,94,-18</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>94 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95,-37,95,-15</points>
<connection>
<GID>2</GID>
<name>IN_B_1</name></connection>
<connection>
<GID>1</GID>
<name>OUT_1</name></connection>
<intersection>-23 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>89.5,-23,95,-23</points>
<connection>
<GID>13</GID>
<name>IN_0</name></connection>
<intersection>95 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96,-37,96,-15</points>
<connection>
<GID>2</GID>
<name>IN_B_0</name></connection>
<connection>
<GID>1</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96.5,-7,96.5,0.5</points>
<connection>
<GID>1</GID>
<name>IN_B_3</name></connection>
<intersection>0.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>97,0.5,97,7.5</points>
<connection>
<GID>3</GID>
<name>OUT_0</name></connection>
<intersection>0.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>96.5,0.5,97,0.5</points>
<intersection>96.5 0</intersection>
<intersection>97 1</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97.5,-7,97.5,0.5</points>
<connection>
<GID>1</GID>
<name>IN_B_2</name></connection>
<intersection>0.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>99,0.5,99,7.5</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>0.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>97.5,0.5,99,0.5</points>
<intersection>97.5 0</intersection>
<intersection>99 1</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>98.5,-7,98.5,0</points>
<connection>
<GID>1</GID>
<name>IN_B_1</name></connection>
<intersection>0 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>101,0,101,7.5</points>
<connection>
<GID>5</GID>
<name>OUT_0</name></connection>
<intersection>0 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>98.5,0,101,0</points>
<intersection>98.5 0</intersection>
<intersection>101 1</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99.5,-7,99.5,-1</points>
<connection>
<GID>1</GID>
<name>IN_B_0</name></connection>
<intersection>-1 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>103,-1,103,7.5</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>-1 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>99.5,-1,103,-1</points>
<intersection>99.5 0</intersection>
<intersection>103 1</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>92.5,-7,92.5,0.5</points>
<connection>
<GID>1</GID>
<name>IN_0</name></connection>
<intersection>0.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>93.5,0.5,93.5,7.5</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>0.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>92.5,0.5,93.5,0.5</points>
<intersection>92.5 0</intersection>
<intersection>93.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91.5,-7,91.5,7.5</points>
<connection>
<GID>1</GID>
<name>IN_1</name></connection>
<connection>
<GID>9</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-7,90.5,0.5</points>
<connection>
<GID>1</GID>
<name>IN_2</name></connection>
<intersection>0.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>89.5,0.5,89.5,7.5</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>0.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>89.5,0.5,90.5,0.5</points>
<intersection>89.5 1</intersection>
<intersection>90.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-7,89.5,-1</points>
<connection>
<GID>1</GID>
<name>IN_3</name></connection>
<intersection>-1 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>87.5,-1,87.5,7.5</points>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection>
<intersection>-1 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>87.5,-1,89.5,-1</points>
<intersection>87.5 1</intersection>
<intersection>89.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83.5,-14,83.5,-10</points>
<intersection>-14 1</intersection>
<intersection>-10 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80.5,-14,83.5,-14</points>
<connection>
<GID>11</GID>
<name>IN_2</name></connection>
<intersection>83.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>83.5,-10,86.5,-10</points>
<connection>
<GID>1</GID>
<name>carry_out</name></connection>
<intersection>83.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82,-17,82,-16</points>
<intersection>-17 1</intersection>
<intersection>-16 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>82,-17,83.5,-17</points>
<connection>
<GID>12</GID>
<name>OUT</name></connection>
<intersection>82 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>80.5,-16,82,-16</points>
<connection>
<GID>11</GID>
<name>IN_1</name></connection>
<intersection>82 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82,-22,82,-18</points>
<intersection>-22 1</intersection>
<intersection>-18 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>82,-22,83.5,-22</points>
<connection>
<GID>13</GID>
<name>OUT</name></connection>
<intersection>82 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>80.5,-18,82,-18</points>
<connection>
<GID>11</GID>
<name>IN_0</name></connection>
<intersection>82 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>86,-35,89,-35</points>
<intersection>86 4</intersection>
<intersection>89 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>89,-37,89,-35</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>-35 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>86,-37,86,-35</points>
<connection>
<GID>2</GID>
<name>IN_3</name></connection>
<intersection>-35 1</intersection></vsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-46,89.5,-45</points>
<connection>
<GID>2</GID>
<name>OUT_3</name></connection>
<intersection>-46 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>86,-48.5,86,-46</points>
<connection>
<GID>17</GID>
<name>N_in3</name></connection>
<intersection>-46 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>86,-46,89.5,-46</points>
<intersection>86 1</intersection>
<intersection>89.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-46.5,90.5,-45</points>
<connection>
<GID>2</GID>
<name>OUT_2</name></connection>
<intersection>-46.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>88.5,-48.5,88.5,-46.5</points>
<connection>
<GID>16</GID>
<name>N_in3</name></connection>
<intersection>-46.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>88.5,-46.5,90.5,-46.5</points>
<intersection>88.5 1</intersection>
<intersection>90.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91.5,-46.5,91.5,-45</points>
<connection>
<GID>2</GID>
<name>OUT_1</name></connection>
<intersection>-46.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>91,-48.5,91,-46.5</points>
<connection>
<GID>15</GID>
<name>N_in3</name></connection>
<intersection>-46.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>91,-46.5,91.5,-46.5</points>
<intersection>91 1</intersection>
<intersection>91.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>92.5,-46.5,92.5,-45</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>-46.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>93.5,-48.5,93.5,-46.5</points>
<connection>
<GID>14</GID>
<name>N_in3</name></connection>
<intersection>-46.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>92.5,-46.5,93.5,-46.5</points>
<intersection>92.5 0</intersection>
<intersection>93.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,-35.5,52.5,-13.5</points>
<connection>
<GID>21</GID>
<name>IN_B_3</name></connection>
<connection>
<GID>20</GID>
<name>OUT_3</name></connection>
<intersection>-19.5 7</intersection>
<intersection>-14.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>49,-14.5,52.5,-14.5</points>
<connection>
<GID>31</GID>
<name>IN_1</name></connection>
<intersection>52.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>49,-19.5,52.5,-19.5</points>
<connection>
<GID>32</GID>
<name>IN_1</name></connection>
<intersection>52.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53.5,-35.5,53.5,-13.5</points>
<connection>
<GID>21</GID>
<name>IN_B_2</name></connection>
<connection>
<GID>20</GID>
<name>OUT_2</name></connection>
<intersection>-16.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>49,-16.5,53.5,-16.5</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>53.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-35.5,54.5,-13.5</points>
<connection>
<GID>21</GID>
<name>IN_B_1</name></connection>
<connection>
<GID>20</GID>
<name>OUT_1</name></connection>
<intersection>-21.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>49,-21.5,54.5,-21.5</points>
<connection>
<GID>32</GID>
<name>IN_0</name></connection>
<intersection>54.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55.5,-35.5,55.5,-13.5</points>
<connection>
<GID>21</GID>
<name>IN_B_0</name></connection>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-5.5,56,2</points>
<connection>
<GID>20</GID>
<name>IN_B_3</name></connection>
<intersection>2 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>56.5,2,56.5,9</points>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection>
<intersection>2 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>56,2,56.5,2</points>
<intersection>56 0</intersection>
<intersection>56.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-5.5,57,2</points>
<connection>
<GID>20</GID>
<name>IN_B_2</name></connection>
<intersection>2 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>58.5,2,58.5,9</points>
<connection>
<GID>23</GID>
<name>OUT_0</name></connection>
<intersection>2 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>57,2,58.5,2</points>
<intersection>57 0</intersection>
<intersection>58.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58,-5.5,58,1.5</points>
<connection>
<GID>20</GID>
<name>IN_B_1</name></connection>
<intersection>1.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>60.5,1.5,60.5,9</points>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection>
<intersection>1.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>58,1.5,60.5,1.5</points>
<intersection>58 0</intersection>
<intersection>60.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59,-5.5,59,0.5</points>
<connection>
<GID>20</GID>
<name>IN_B_0</name></connection>
<intersection>0.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>62.5,0.5,62.5,9</points>
<connection>
<GID>25</GID>
<name>OUT_0</name></connection>
<intersection>0.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>59,0.5,62.5,0.5</points>
<intersection>59 0</intersection>
<intersection>62.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,-5.5,52,2</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>2 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>53,2,53,9</points>
<connection>
<GID>29</GID>
<name>OUT_0</name></connection>
<intersection>2 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>52,2,53,2</points>
<intersection>52 0</intersection>
<intersection>53 1</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51,-5.5,51,9</points>
<connection>
<GID>20</GID>
<name>IN_1</name></connection>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50,-5.5,50,2</points>
<connection>
<GID>20</GID>
<name>IN_2</name></connection>
<intersection>2 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>49,2,49,9</points>
<connection>
<GID>27</GID>
<name>OUT_0</name></connection>
<intersection>2 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>49,2,50,2</points>
<intersection>49 1</intersection>
<intersection>50 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,-5.5,49,0.5</points>
<connection>
<GID>20</GID>
<name>IN_3</name></connection>
<intersection>0.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>47,0.5,47,9</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<intersection>0.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>47,0.5,49,0.5</points>
<intersection>47 1</intersection>
<intersection>49 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43,-12.5,43,-8.5</points>
<intersection>-12.5 1</intersection>
<intersection>-8.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40,-12.5,43,-12.5</points>
<connection>
<GID>30</GID>
<name>IN_2</name></connection>
<intersection>43 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>43,-8.5,46,-8.5</points>
<connection>
<GID>20</GID>
<name>carry_out</name></connection>
<intersection>43 0</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41.5,-15.5,41.5,-14.5</points>
<intersection>-15.5 1</intersection>
<intersection>-14.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41.5,-15.5,43,-15.5</points>
<connection>
<GID>31</GID>
<name>OUT</name></connection>
<intersection>41.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>40,-14.5,41.5,-14.5</points>
<connection>
<GID>30</GID>
<name>IN_1</name></connection>
<intersection>41.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41.5,-20.5,41.5,-16.5</points>
<intersection>-20.5 1</intersection>
<intersection>-16.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41.5,-20.5,43,-20.5</points>
<connection>
<GID>32</GID>
<name>OUT</name></connection>
<intersection>41.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>40,-16.5,41.5,-16.5</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>41.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,-29.5,47.5,-29.5</points>
<intersection>34 3</intersection>
<intersection>46.5 9</intersection>
<intersection>47.5 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>34,-46.5,34,-14.5</points>
<connection>
<GID>30</GID>
<name>OUT</name></connection>
<intersection>-46.5 7</intersection>
<intersection>-29.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>47.5,-35.5,47.5,-29.5</points>
<connection>
<GID>21</GID>
<name>IN_1</name></connection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>34,-46.5,39.5,-46.5</points>
<connection>
<GID>37</GID>
<name>N_in3</name></connection>
<intersection>34 3</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>46.5,-35.5,46.5,-29.5</points>
<connection>
<GID>21</GID>
<name>IN_2</name></connection>
<intersection>-29.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-33.5,48.5,-33.5</points>
<intersection>45.5 4</intersection>
<intersection>48.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>48.5,-35.5,48.5,-33.5</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<intersection>-33.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>45.5,-35.5,45.5,-33.5</points>
<connection>
<GID>21</GID>
<name>IN_3</name></connection>
<intersection>-33.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,-44.5,49,-43.5</points>
<connection>
<GID>21</GID>
<name>OUT_3</name></connection>
<intersection>-44.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>45.5,-47,45.5,-44.5</points>
<connection>
<GID>36</GID>
<name>N_in3</name></connection>
<intersection>-44.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>45.5,-44.5,49,-44.5</points>
<intersection>45.5 1</intersection>
<intersection>49 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50,-45,50,-43.5</points>
<connection>
<GID>21</GID>
<name>OUT_2</name></connection>
<intersection>-45 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>48,-47,48,-45</points>
<connection>
<GID>35</GID>
<name>N_in3</name></connection>
<intersection>-45 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>48,-45,50,-45</points>
<intersection>48 1</intersection>
<intersection>50 0</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51,-45,51,-43.5</points>
<connection>
<GID>21</GID>
<name>OUT_1</name></connection>
<intersection>-45 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>50.5,-47,50.5,-45</points>
<connection>
<GID>34</GID>
<name>N_in3</name></connection>
<intersection>-45 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>50.5,-45,51,-45</points>
<intersection>50.5 1</intersection>
<intersection>51 0</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,-45,52,-43.5</points>
<connection>
<GID>21</GID>
<name>OUT_0</name></connection>
<intersection>-45 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>53,-47,53,-45</points>
<connection>
<GID>33</GID>
<name>N_in3</name></connection>
<intersection>-45 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>52,-45,53,-45</points>
<intersection>52 0</intersection>
<intersection>53 1</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-33,88,-33</points>
<intersection>73.5 2</intersection>
<intersection>87 6</intersection>
<intersection>88 7</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>73.5,-33,73.5,-16</points>
<intersection>-33 1</intersection>
<intersection>-16 5</intersection></vsegment>
<vsegment>
<ID>3</ID>
<points>68,-16,68,-8.5</points>
<intersection>-16 5</intersection>
<intersection>-8.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>62,-8.5,68,-8.5</points>
<connection>
<GID>20</GID>
<name>carry_in</name></connection>
<intersection>68 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>68,-16,74.5,-16</points>
<connection>
<GID>11</GID>
<name>OUT</name></connection>
<intersection>68 3</intersection>
<intersection>73.5 2</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>87,-37,87,-33</points>
<connection>
<GID>2</GID>
<name>IN_2</name></connection>
<intersection>-33 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>88,-37,88,-33</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>-33 1</intersection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 1>
<page 2>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 2>
<page 3>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 3>
<page 4>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 4>
<page 5>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 5>
<page 6>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 6>
<page 7>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 7>
<page 8>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 8>
<page 9>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 9></circuit>