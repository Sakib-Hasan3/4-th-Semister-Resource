<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-23.0667,0.7,116.333,-69.5</PageViewport>
<gate>
<ID>2</ID>
<type>AA_AND2</type>
<position>19,-15</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_INVERTER</type>
<position>19,-9.5</position>
<input>
<ID>IN_0</ID>2 </input>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6</ID>
<type>AE_OR2</type>
<position>19,-22</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_INVERTER</type>
<position>18,-34.5</position>
<input>
<ID>IN_0</ID>4 </input>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_INVERTER</type>
<position>29,-22</position>
<input>
<ID>IN_0</ID>7 </input>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>12</ID>
<type>AE_OR2</type>
<position>38,-16</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_AND2</type>
<position>38,-22.5</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>4 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_AND2</type>
<position>38,-33.5</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>8 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_AND2</type>
<position>38,-40.5</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>4 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>20</ID>
<type>AE_OR2</type>
<position>50,-41.5</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>22</ID>
<type>AE_OR2</type>
<position>50,-25.5</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_TOGGLE</type>
<position>1,-13.5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_TOGGLE</type>
<position>1,-27</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_TOGGLE</type>
<position>1,-19</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>30</ID>
<type>AA_TOGGLE</type>
<position>1.5,-44</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>32</ID>
<type>GA_LED</type>
<position>63,-7.5</position>
<input>
<ID>N_in0</ID>1 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>GA_LED</type>
<position>63,-16.5</position>
<input>
<ID>N_in0</ID>13 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>36</ID>
<type>GA_LED</type>
<position>63,-25.5</position>
<input>
<ID>N_in0</ID>14 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>38</ID>
<type>GA_LED</type>
<position>63,-36.5</position>
<input>
<ID>N_in0</ID>15 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>40</ID>
<type>AA_LABEL</type>
<position>-6,-44</position>
<gparam>LABEL_TEXT A0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>41</ID>
<type>AA_LABEL</type>
<position>67,-36.5</position>
<gparam>LABEL_TEXT E0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>42</ID>
<type>AA_LABEL</type>
<position>67,-25</position>
<gparam>LABEL_TEXT E1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>43</ID>
<type>AA_LABEL</type>
<position>67.5,-16.5</position>
<gparam>LABEL_TEXT E2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>44</ID>
<type>AA_LABEL</type>
<position>67.5,-7.5</position>
<gparam>LABEL_TEXT E3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>45</ID>
<type>AA_LABEL</type>
<position>-6,-27</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>46</ID>
<type>AA_LABEL</type>
<position>-5.5,-19</position>
<gparam>LABEL_TEXT A2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>47</ID>
<type>AA_LABEL</type>
<position>-5.5,-13</position>
<gparam>LABEL_TEXT A3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42,-9.5,42,-7.5</points>
<intersection>-9.5 2</intersection>
<intersection>-7.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>42,-7.5,62,-7.5</points>
<connection>
<GID>32</GID>
<name>N_in0</name></connection>
<intersection>42 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22,-9.5,42,-9.5</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>42 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3,-13.5,16,-13.5</points>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection>
<intersection>9 4</intersection>
<intersection>13.5 6</intersection>
<intersection>16 11</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>9,-13.5,9,-9.5</points>
<intersection>-13.5 1</intersection>
<intersection>-9.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>9,-9.5,16,-9.5</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>9 4</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>13.5,-21,13.5,-13.5</points>
<intersection>-21 7</intersection>
<intersection>-13.5 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>13.5,-21,16,-21</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>13.5 6</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>16,-14,16,-13.5</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>-13.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,-23,11,-16</points>
<intersection>-23 3</intersection>
<intersection>-19 2</intersection>
<intersection>-16 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>11,-16,16,-16</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>11 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>3,-19,11,-19</points>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection>
<intersection>11 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>11,-23,16,-23</points>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<intersection>11 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3,-27,32,-27</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<intersection>8.5 9</intersection>
<intersection>32 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>32,-27,32,-23.5</points>
<intersection>-27 1</intersection>
<intersection>-23.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>32,-23.5,35,-23.5</points>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<intersection>32 3</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>8.5,-41.5,8.5,-27</points>
<intersection>-41.5 10</intersection>
<intersection>-34.5 12</intersection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>8.5,-41.5,35,-41.5</points>
<connection>
<GID>18</GID>
<name>IN_1</name></connection>
<intersection>8.5 9</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>8.5,-34.5,15,-34.5</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>8.5 9</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22,-15,35,-15</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<connection>
<GID>2</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33.5,-22,33.5,-17</points>
<intersection>-22 2</intersection>
<intersection>-21.5 3</intersection>
<intersection>-17 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33.5,-17,35,-17</points>
<connection>
<GID>12</GID>
<name>IN_1</name></connection>
<intersection>33.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32,-22,33.5,-22</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>33.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>33.5,-21.5,35,-21.5</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>33.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22,-22,26,-22</points>
<connection>
<GID>6</GID>
<name>OUT</name></connection>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>24.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>24.5,-39.5,24.5,-22</points>
<intersection>-39.5 6</intersection>
<intersection>-32.5 4</intersection>
<intersection>-22 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>24.5,-32.5,35,-32.5</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>24.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>24.5,-39.5,35,-39.5</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>24.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>21,-34.5,35,-34.5</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,-40.5,47,-40.5</points>
<connection>
<GID>18</GID>
<name>OUT</name></connection>
<connection>
<GID>20</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3.5,-44,47,-44</points>
<connection>
<GID>30</GID>
<name>OUT_0</name></connection>
<intersection>47 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>47,-44,47,-42.5</points>
<connection>
<GID>20</GID>
<name>IN_1</name></connection>
<intersection>-44 1</intersection></vsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44,-33.5,44,-26.5</points>
<intersection>-33.5 2</intersection>
<intersection>-26.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44,-26.5,47,-26.5</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<intersection>44 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>41,-33.5,44,-33.5</points>
<connection>
<GID>16</GID>
<name>OUT</name></connection>
<intersection>44 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44,-24.5,44,-22.5</points>
<intersection>-24.5 1</intersection>
<intersection>-22.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44,-24.5,47,-24.5</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>44 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>41,-22.5,44,-22.5</points>
<connection>
<GID>14</GID>
<name>OUT</name></connection>
<intersection>44 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51.5,-16.5,51.5,-16</points>
<intersection>-16.5 1</intersection>
<intersection>-16 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51.5,-16.5,62,-16.5</points>
<connection>
<GID>34</GID>
<name>N_in0</name></connection>
<intersection>51.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>41,-16,51.5,-16</points>
<connection>
<GID>12</GID>
<name>OUT</name></connection>
<intersection>51.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-25.5,62,-25.5</points>
<connection>
<GID>36</GID>
<name>N_in0</name></connection>
<connection>
<GID>22</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57.5,-41.5,57.5,-36.5</points>
<intersection>-41.5 2</intersection>
<intersection>-36.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>57.5,-36.5,62,-36.5</points>
<connection>
<GID>38</GID>
<name>N_in0</name></connection>
<intersection>57.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>53,-41.5,57.5,-41.5</points>
<connection>
<GID>20</GID>
<name>OUT</name></connection>
<intersection>57.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 1>
<page 2>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 2>
<page 3>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 3>
<page 4>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 4>
<page 5>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 5>
<page 6>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 6>
<page 7>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 7>
<page 8>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 8>
<page 9>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 9></circuit>