<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>0,0,139.4,-70.2</PageViewport>
<gate>
<ID>2</ID>
<type>AA_TOGGLE</type>
<position>20,-7</position>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>25.5,-7</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>5</ID>
<type>AA_TOGGLE</type>
<position>38.5,-7</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>44.5,-7</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_INVERTER</type>
<position>29.5,-19.5</position>
<input>
<ID>IN_0</ID>1 </input>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>10</ID>
<type>GA_LED</type>
<position>61.5,-19</position>
<input>
<ID>N_in0</ID>2 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>AA_AND2</type>
<position>42,-27</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>1 </input>
<output>
<ID>OUT</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>13</ID>
<type>AA_AND2</type>
<position>42,-32</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>15</ID>
<type>AE_OR2</type>
<position>50,-29</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>4 </input>
<output>
<ID>OUT</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>16</ID>
<type>GA_LED</type>
<position>61.5,-29</position>
<input>
<ID>N_in0</ID>5 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>19</ID>
<type>AA_INVERTER</type>
<position>41,-19.5</position>
<input>
<ID>IN_0</ID>6 </input>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_INVERTER</type>
<position>24.5,-19.5</position>
<input>
<ID>IN_0</ID>8 </input>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_AND2</type>
<position>42,-41</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_AND2</type>
<position>42,-46</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>12 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_AND3</type>
<position>42,-52</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>7 </input>
<input>
<ID>IN_2</ID>2 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>28</ID>
<type>AE_OR3</type>
<position>52.5,-46</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>10 </input>
<input>
<ID>IN_2</ID>11 </input>
<output>
<ID>OUT</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>29</ID>
<type>GA_LED</type>
<position>62,-46</position>
<input>
<ID>N_in0</ID>13 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>31</ID>
<type>AA_AND2</type>
<position>42,-61</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>33</ID>
<type>AA_AND2</type>
<position>42,-65.5</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>1 </input>
<output>
<ID>OUT</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>35</ID>
<type>AE_OR3</type>
<position>52,-63</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>15 </input>
<input>
<ID>IN_2</ID>16 </input>
<output>
<ID>OUT</ID>17 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>36</ID>
<type>GA_LED</type>
<position>62,-62.5</position>
<input>
<ID>N_in0</ID>17 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36.5,-28,36.5,-11</points>
<intersection>-28 3</intersection>
<intersection>-11 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>31.5,-28,39,-28</points>
<connection>
<GID>12</GID>
<name>IN_1</name></connection>
<intersection>31.5 8</intersection>
<intersection>36.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>29.5,-11,44.5,-11</points>
<intersection>29.5 7</intersection>
<intersection>36.5 0</intersection>
<intersection>44.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>44.5,-11,44.5,-9</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>-11 4</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>29.5,-16.5,29.5,-11</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>-11 4</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>31.5,-45,31.5,-28</points>
<intersection>-45 9</intersection>
<intersection>-28 3</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>31.5,-45,39,-45</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>31.5 8</intersection>
<intersection>38 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>38,-66.5,38,-45</points>
<intersection>-66.5 11</intersection>
<intersection>-45 9</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>38,-66.5,39,-66.5</points>
<connection>
<GID>33</GID>
<name>IN_1</name></connection>
<intersection>38 10</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-33,32.5,-19</points>
<intersection>-33 5</intersection>
<intersection>-22.5 4</intersection>
<intersection>-19 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32.5,-19,60.5,-19</points>
<connection>
<GID>10</GID>
<name>N_in0</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>29.5,-22.5,32.5,-22.5</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>30.5,-33,39,-33</points>
<connection>
<GID>13</GID>
<name>IN_1</name></connection>
<intersection>30.5 6</intersection>
<intersection>32.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>30.5,-54,30.5,-33</points>
<intersection>-54 7</intersection>
<intersection>-33 5</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>30.5,-54,39,-54</points>
<connection>
<GID>26</GID>
<name>IN_2</name></connection>
<intersection>30.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46,-28,46,-27</points>
<intersection>-28 1</intersection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46,-28,47,-28</points>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<intersection>46 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>45,-27,46,-27</points>
<connection>
<GID>12</GID>
<name>OUT</name></connection>
<intersection>46 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46,-32,46,-30</points>
<intersection>-32 2</intersection>
<intersection>-30 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46,-30,47,-30</points>
<connection>
<GID>15</GID>
<name>IN_1</name></connection>
<intersection>46 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>45,-32,46,-32</points>
<connection>
<GID>13</GID>
<name>OUT</name></connection>
<intersection>46 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-29,60.5,-29</points>
<connection>
<GID>16</GID>
<name>N_in0</name></connection>
<connection>
<GID>15</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,-26,38.5,-9</points>
<connection>
<GID>5</GID>
<name>OUT_0</name></connection>
<intersection>-26 1</intersection>
<intersection>-16.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34.5,-26,39,-26</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>34.5 3</intersection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>38.5,-16.5,41,-16.5</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<intersection>38.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>34.5,-42,34.5,-26</points>
<intersection>-42 4</intersection>
<intersection>-26 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>33.5,-42,39,-42</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<intersection>33.5 5</intersection>
<intersection>34.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>33.5,-62,33.5,-42</points>
<intersection>-62 6</intersection>
<intersection>-42 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>33.5,-62,39,-62</points>
<connection>
<GID>31</GID>
<name>IN_1</name></connection>
<intersection>33.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33.5,-31,33.5,-22.5</points>
<intersection>-31 1</intersection>
<intersection>-22.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33.5,-31,39,-31</points>
<connection>
<GID>13</GID>
<name>IN_0</name></connection>
<intersection>33.5 0</intersection>
<intersection>36.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>33.5,-22.5,41,-22.5</points>
<connection>
<GID>19</GID>
<name>OUT_0</name></connection>
<intersection>33.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>36.5,-52,36.5,-31</points>
<intersection>-52 4</intersection>
<intersection>-31 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>36.5,-52,39,-52</points>
<connection>
<GID>26</GID>
<name>IN_1</name></connection>
<intersection>36.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-50,22.5,-12.5</points>
<intersection>-50 3</intersection>
<intersection>-16.5 4</intersection>
<intersection>-12.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>25.5,-12.5,25.5,-9</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>-12.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>22.5,-12.5,25.5,-12.5</points>
<intersection>22.5 0</intersection>
<intersection>25.5 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>22.5,-50,39,-50</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>22.5 0</intersection>
<intersection>35 5</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>22.5,-16.5,24.5,-16.5</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>22.5 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>35,-60,35,-50</points>
<intersection>-60 6</intersection>
<intersection>-50 3</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>35,-60,39,-60</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>35 5</intersection>
<intersection>37 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>37,-64.5,37,-60</points>
<intersection>-64.5 8</intersection>
<intersection>-60 6</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>37,-64.5,39,-64.5</points>
<connection>
<GID>33</GID>
<name>IN_0</name></connection>
<intersection>37 7</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,-44,47,-41</points>
<intersection>-44 1</intersection>
<intersection>-41 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,-44,49.5,-44</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<intersection>47 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>45,-41,47,-41</points>
<connection>
<GID>22</GID>
<name>OUT</name></connection>
<intersection>47 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-46,49.5,-46</points>
<connection>
<GID>28</GID>
<name>IN_1</name></connection>
<connection>
<GID>24</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,-52,47,-48</points>
<intersection>-52 2</intersection>
<intersection>-48 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,-48,49.5,-48</points>
<connection>
<GID>28</GID>
<name>IN_2</name></connection>
<intersection>47 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>45,-52,47,-52</points>
<connection>
<GID>26</GID>
<name>OUT</name></connection>
<intersection>47 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-40,24.5,-22.5</points>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<intersection>-40 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24.5,-40,39,-40</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>24.5 0</intersection>
<intersection>38 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>38,-47,38,-40</points>
<intersection>-47 3</intersection>
<intersection>-40 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>38,-47,39,-47</points>
<connection>
<GID>24</GID>
<name>IN_1</name></connection>
<intersection>38 2</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55.5,-46,61,-46</points>
<connection>
<GID>29</GID>
<name>N_in0</name></connection>
<connection>
<GID>28</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-61,49,-61</points>
<connection>
<GID>35</GID>
<name>IN_0</name></connection>
<connection>
<GID>31</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,-65.5,47,-63</points>
<intersection>-65.5 2</intersection>
<intersection>-63 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,-63,49,-63</points>
<connection>
<GID>35</GID>
<name>IN_1</name></connection>
<intersection>47 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>45,-65.5,47,-65.5</points>
<connection>
<GID>33</GID>
<name>OUT</name></connection>
<intersection>47 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20,-68,20,-9</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>-68 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20,-68,49,-68</points>
<intersection>20 0</intersection>
<intersection>49 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>49,-68,49,-65</points>
<connection>
<GID>35</GID>
<name>IN_2</name></connection>
<intersection>-68 1</intersection></vsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58,-63,58,-62.5</points>
<intersection>-63 2</intersection>
<intersection>-62.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58,-62.5,61,-62.5</points>
<connection>
<GID>36</GID>
<name>N_in0</name></connection>
<intersection>58 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>55,-63,58,-63</points>
<connection>
<GID>35</GID>
<name>OUT</name></connection>
<intersection>58 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 1>
<page 2>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 2>
<page 3>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 3>
<page 4>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 4>
<page 5>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 5>
<page 6>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 6>
<page 7>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 7>
<page 8>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 8>
<page 9>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 9></circuit>