<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-0.997949,16.8786,153.716,-61.0335</PageViewport>
<gate>
<ID>2</ID>
<type>AE_FULLADDER_4BIT</type>
<position>65.5,-18</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>10 </input>
<input>
<ID>IN_2</ID>11 </input>
<input>
<ID>IN_3</ID>12 </input>
<input>
<ID>IN_B_0</ID>8 </input>
<input>
<ID>IN_B_1</ID>7 </input>
<input>
<ID>IN_B_2</ID>6 </input>
<input>
<ID>IN_B_3</ID>5 </input>
<output>
<ID>OUT_0</ID>4 </output>
<output>
<ID>OUT_1</ID>3 </output>
<output>
<ID>OUT_2</ID>2 </output>
<output>
<ID>OUT_3</ID>1 </output>
<output>
<ID>carry_out</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>4</ID>
<type>AE_FULLADDER_4BIT</type>
<position>62,-48</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>16 </input>
<input>
<ID>IN_2</ID>16 </input>
<input>
<ID>IN_3</ID>17 </input>
<input>
<ID>IN_B_0</ID>4 </input>
<input>
<ID>IN_B_1</ID>3 </input>
<input>
<ID>IN_B_2</ID>2 </input>
<input>
<ID>IN_B_3</ID>1 </input>
<output>
<ID>OUT_0</ID>21 </output>
<output>
<ID>OUT_1</ID>20 </output>
<output>
<ID>OUT_2</ID>19 </output>
<output>
<ID>OUT_3</ID>18 </output>
<output>
<ID>carry_out</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>68,2.5</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>7</ID>
<type>AA_TOGGLE</type>
<position>70,2.5</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_TOGGLE</type>
<position>72,2.5</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>9</ID>
<type>AA_TOGGLE</type>
<position>74,2.5</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_TOGGLE</type>
<position>58.5,2.5</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>15</ID>
<type>AA_TOGGLE</type>
<position>60.5,2.5</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_TOGGLE</type>
<position>62.5,2.5</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>17</ID>
<type>AA_TOGGLE</type>
<position>64.5,2.5</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>19</ID>
<type>AE_OR3</type>
<position>48.5,-23</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>14 </input>
<input>
<ID>IN_2</ID>13 </input>
<output>
<ID>OUT</ID>16 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>21</ID>
<type>AA_AND2</type>
<position>57.5,-24</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>1 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>23</ID>
<type>AA_AND2</type>
<position>57.5,-29</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>1 </input>
<output>
<ID>OUT</ID>15 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>25</ID>
<type>GA_LED</type>
<position>64.5,-56.5</position>
<input>
<ID>N_in3</ID>21 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>27</ID>
<type>GA_LED</type>
<position>62,-56.5</position>
<input>
<ID>N_in3</ID>20 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>29</ID>
<type>GA_LED</type>
<position>59.5,-56.5</position>
<input>
<ID>N_in3</ID>19 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>31</ID>
<type>GA_LED</type>
<position>57,-56.5</position>
<input>
<ID>N_in3</ID>18 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>33</ID>
<type>GA_LED</type>
<position>51,-56</position>
<input>
<ID>N_in3</ID>16 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>35</ID>
<type>GA_LED</type>
<position>50.5,-46.5</position>
<input>
<ID>N_in1</ID>22 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64,-44,64,-22</points>
<connection>
<GID>2</GID>
<name>OUT_3</name></connection>
<connection>
<GID>4</GID>
<name>IN_B_3</name></connection>
<intersection>-28 7</intersection>
<intersection>-23 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>60.5,-23,64,-23</points>
<connection>
<GID>21</GID>
<name>IN_1</name></connection>
<intersection>64 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>60.5,-28,64,-28</points>
<connection>
<GID>23</GID>
<name>IN_1</name></connection>
<intersection>64 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65,-44,65,-22</points>
<connection>
<GID>2</GID>
<name>OUT_2</name></connection>
<connection>
<GID>4</GID>
<name>IN_B_2</name></connection>
<intersection>-25 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>60.5,-25,65,-25</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<intersection>65 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66,-44,66,-22</points>
<connection>
<GID>2</GID>
<name>OUT_1</name></connection>
<connection>
<GID>4</GID>
<name>IN_B_1</name></connection>
<intersection>-30 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>60.5,-30,66,-30</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<intersection>66 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67,-44,67,-22</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<connection>
<GID>4</GID>
<name>IN_B_0</name></connection></vsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67.5,-14,67.5,-6.5</points>
<connection>
<GID>2</GID>
<name>IN_B_3</name></connection>
<intersection>-6.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>68,-6.5,68,0.5</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>-6.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>67.5,-6.5,68,-6.5</points>
<intersection>67.5 0</intersection>
<intersection>68 1</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68.5,-14,68.5,-6.5</points>
<connection>
<GID>2</GID>
<name>IN_B_2</name></connection>
<intersection>-6.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>70,-6.5,70,0.5</points>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection>
<intersection>-6.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>68.5,-6.5,70,-6.5</points>
<intersection>68.5 0</intersection>
<intersection>70 1</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69.5,-14,69.5,-7</points>
<connection>
<GID>2</GID>
<name>IN_B_1</name></connection>
<intersection>-7 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>72,-7,72,0.5</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>-7 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>69.5,-7,72,-7</points>
<intersection>69.5 0</intersection>
<intersection>72 1</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70.5,-14,70.5,-8</points>
<connection>
<GID>2</GID>
<name>IN_B_0</name></connection>
<intersection>-8 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>74,-8,74,0.5</points>
<connection>
<GID>9</GID>
<name>OUT_0</name></connection>
<intersection>-8 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>70.5,-8,74,-8</points>
<intersection>70.5 0</intersection>
<intersection>74 1</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63.5,-14,63.5,-6.5</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>-6.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>64.5,-6.5,64.5,0.5</points>
<connection>
<GID>17</GID>
<name>OUT_0</name></connection>
<intersection>-6.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>63.5,-6.5,64.5,-6.5</points>
<intersection>63.5 0</intersection>
<intersection>64.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62.5,-14,62.5,0.5</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61.5,-14,61.5,-6.5</points>
<connection>
<GID>2</GID>
<name>IN_2</name></connection>
<intersection>-6.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>60.5,-6.5,60.5,0.5</points>
<connection>
<GID>15</GID>
<name>OUT_0</name></connection>
<intersection>-6.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>60.5,-6.5,61.5,-6.5</points>
<intersection>60.5 1</intersection>
<intersection>61.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,-14,60.5,-8</points>
<connection>
<GID>2</GID>
<name>IN_3</name></connection>
<intersection>-8 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>58.5,-8,58.5,0.5</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>-8 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>58.5,-8,60.5,-8</points>
<intersection>58.5 1</intersection>
<intersection>60.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-21,54.5,-17</points>
<intersection>-21 1</intersection>
<intersection>-17 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51.5,-21,54.5,-21</points>
<connection>
<GID>19</GID>
<name>IN_2</name></connection>
<intersection>54.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>54.5,-17,57.5,-17</points>
<connection>
<GID>2</GID>
<name>carry_out</name></connection>
<intersection>54.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,-24,53,-23</points>
<intersection>-24 1</intersection>
<intersection>-23 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53,-24,54.5,-24</points>
<connection>
<GID>21</GID>
<name>OUT</name></connection>
<intersection>53 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>51.5,-23,53,-23</points>
<connection>
<GID>19</GID>
<name>IN_1</name></connection>
<intersection>53 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,-29,53,-25</points>
<intersection>-29 1</intersection>
<intersection>-25 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53,-29,54.5,-29</points>
<connection>
<GID>23</GID>
<name>OUT</name></connection>
<intersection>53 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>51.5,-25,53,-25</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<intersection>53 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-38,59,-38</points>
<intersection>45.5 3</intersection>
<intersection>58 9</intersection>
<intersection>59 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>45.5,-55,45.5,-23</points>
<connection>
<GID>19</GID>
<name>OUT</name></connection>
<intersection>-55 7</intersection>
<intersection>-38 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>59,-44,59,-38</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<intersection>-38 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>45.5,-55,51,-55</points>
<connection>
<GID>33</GID>
<name>N_in3</name></connection>
<intersection>45.5 3</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>58,-44,58,-38</points>
<connection>
<GID>4</GID>
<name>IN_2</name></connection>
<intersection>-38 1</intersection></vsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57,-42,60,-42</points>
<intersection>57 4</intersection>
<intersection>60 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>60,-44,60,-42</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>-42 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>57,-44,57,-42</points>
<connection>
<GID>4</GID>
<name>IN_3</name></connection>
<intersection>-42 1</intersection></vsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,-53,60.5,-52</points>
<connection>
<GID>4</GID>
<name>OUT_3</name></connection>
<intersection>-53 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>57,-55.5,57,-53</points>
<connection>
<GID>31</GID>
<name>N_in3</name></connection>
<intersection>-53 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>57,-53,60.5,-53</points>
<intersection>57 1</intersection>
<intersection>60.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61.5,-53.5,61.5,-52</points>
<connection>
<GID>4</GID>
<name>OUT_2</name></connection>
<intersection>-53.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>59.5,-55.5,59.5,-53.5</points>
<connection>
<GID>29</GID>
<name>N_in3</name></connection>
<intersection>-53.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>59.5,-53.5,61.5,-53.5</points>
<intersection>59.5 1</intersection>
<intersection>61.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62.5,-53.5,62.5,-52</points>
<connection>
<GID>4</GID>
<name>OUT_1</name></connection>
<intersection>-53.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>62,-55.5,62,-53.5</points>
<connection>
<GID>27</GID>
<name>N_in3</name></connection>
<intersection>-53.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>62,-53.5,62.5,-53.5</points>
<intersection>62 1</intersection>
<intersection>62.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63.5,-53.5,63.5,-52</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>-53.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>64.5,-55.5,64.5,-53.5</points>
<connection>
<GID>25</GID>
<name>N_in3</name></connection>
<intersection>-53.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>63.5,-53.5,64.5,-53.5</points>
<intersection>63.5 0</intersection>
<intersection>64.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,-47,52.5,-46.5</points>
<intersection>-47 1</intersection>
<intersection>-46.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52.5,-47,54,-47</points>
<connection>
<GID>4</GID>
<name>carry_out</name></connection>
<intersection>52.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>51.5,-46.5,52.5,-46.5</points>
<connection>
<GID>35</GID>
<name>N_in1</name></connection>
<intersection>52.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 1>
<page 2>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 2>
<page 3>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 3>
<page 4>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 4>
<page 5>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 5>
<page 6>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 6>
<page 7>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 7>
<page 8>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 8>
<page 9>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 9></circuit>